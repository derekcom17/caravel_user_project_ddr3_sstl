magic
tech sky130A
magscale 1 2
timestamp 1644908151
<< checkpaint >>
rect -1242 -1244 10278 24764
rect 12190 13340 34566 36732
rect 11454 10724 34566 13340
rect 11454 10180 14142 10724
<< locali >>
rect 22027 32313 23103 32425
rect 22027 29049 23103 29161
rect 22027 25785 23103 25897
rect 1709 23198 1735 23243
rect 22027 22521 23103 22633
rect 441 20345 442 20407
rect 1709 19934 1735 19979
rect 22027 19257 23103 19369
rect 441 17081 442 17143
rect 1709 16670 1735 16715
rect 22027 15993 23103 16105
rect 441 13817 442 13879
rect 1709 13406 1735 13451
rect 22027 12729 23103 12841
rect 10394 11737 10551 11806
rect 11502 11718 11532 11750
rect 12361 11701 12459 11744
rect 441 10553 442 10615
rect 1709 10142 1735 10187
rect 441 7289 442 7351
rect 1709 6878 1735 6923
rect 441 4025 442 4087
<< viali >>
rect 20671 35167 20709 35205
rect 23165 35161 23215 35211
rect 23358 35159 23402 35203
rect 23542 35138 23586 35182
rect 26057 35166 26091 35200
rect 23103 32313 23215 32425
rect 23358 32380 23402 32424
rect 23450 32380 23494 32424
rect 24734 32314 24778 32358
rect 20671 31903 20709 31941
rect 23165 31897 23215 31947
rect 23358 31895 23402 31939
rect 23542 31874 23586 31918
rect 26057 31902 26091 31936
rect 23103 29049 23215 29161
rect 23358 29116 23402 29160
rect 23450 29116 23494 29160
rect 24734 29050 24778 29094
rect 20671 28639 20709 28677
rect 23165 28633 23215 28683
rect 23358 28631 23402 28675
rect 23542 28610 23586 28654
rect 26057 28638 26091 28672
rect 23103 25785 23215 25897
rect 23358 25852 23402 25896
rect 23450 25852 23494 25896
rect 24734 25786 24778 25830
rect 20671 25375 20709 25413
rect 23165 25369 23215 25419
rect 23358 25367 23402 25411
rect 23542 25346 23586 25390
rect 26057 25374 26091 25408
rect 1769 23209 1803 23243
rect 23103 22521 23215 22633
rect 23358 22588 23402 22632
rect 23450 22588 23494 22632
rect 24734 22522 24778 22566
rect 20671 22111 20709 22149
rect 23165 22105 23215 22155
rect 23358 22103 23402 22147
rect 23542 22082 23586 22126
rect 26057 22110 26091 22144
rect 442 20345 504 20407
rect 1769 19945 1803 19979
rect 23103 19257 23215 19369
rect 23358 19324 23402 19368
rect 23450 19324 23494 19368
rect 24734 19258 24778 19302
rect 20671 18847 20709 18885
rect 23165 18841 23215 18891
rect 23358 18839 23402 18883
rect 23542 18818 23586 18862
rect 26057 18846 26091 18880
rect 442 17081 504 17143
rect 1769 16681 1803 16715
rect 23103 15993 23215 16105
rect 23358 16060 23402 16104
rect 23450 16060 23494 16104
rect 24734 15994 24778 16038
rect 20671 15583 20709 15621
rect 23165 15577 23215 15627
rect 23358 15575 23402 15619
rect 23542 15554 23586 15598
rect 26057 15582 26091 15616
rect 442 13817 504 13879
rect 1769 13417 1803 13451
rect 23103 12729 23215 12841
rect 23358 12796 23402 12840
rect 23450 12796 23494 12840
rect 24734 12730 24778 12774
rect 11111 11830 11159 11878
rect 9807 11637 9873 11703
rect 9993 11678 10061 11746
rect 10178 11684 10234 11740
rect 10626 11737 10700 11811
rect 11412 11749 11461 11798
rect 11532 11717 11566 11751
rect 11663 11737 11721 11795
rect 12679 11752 12735 11808
rect 12459 11701 12504 11746
rect 442 10553 504 10615
rect 1769 10153 1803 10187
rect 442 7289 504 7351
rect 1769 6889 1803 6923
rect 442 4025 504 4087
rect 1769 3625 1803 3659
rect 442 761 504 823
<< metal1 >>
rect 23254 35394 23260 35450
rect 23316 35394 23322 35450
rect 23159 35211 23221 35223
rect 20659 35205 23165 35211
rect 20659 35167 20671 35205
rect 20709 35167 23165 35205
rect 20659 35161 23165 35167
rect 23215 35161 23221 35211
rect 23159 35155 23221 35161
rect 23159 35149 23215 35155
rect 23346 35153 23352 35209
rect 23408 35153 23414 35209
rect 23165 35127 23215 35149
rect 23530 35132 23536 35188
rect 23592 35132 23598 35188
rect 23945 35140 23951 35253
rect 24064 35209 24070 35253
rect 24068 35200 24074 35209
rect 26045 35200 26103 35206
rect 24068 35166 26057 35200
rect 26091 35166 26103 35200
rect 24068 35157 24074 35166
rect 26045 35160 26103 35166
rect 24064 35140 24070 35157
rect 23173 35064 23214 35127
rect 23863 35070 23915 35076
rect 23173 35023 23863 35064
rect 23863 35012 23915 35018
rect 23162 34852 23168 34908
rect 23224 34852 23230 34908
rect 22518 32847 22524 32848
rect 22511 32792 22524 32847
rect 22580 32847 22586 32848
rect 22580 32792 23352 32847
rect 22511 32791 23352 32792
rect 23408 32791 23415 32847
rect 23162 32678 23168 32734
rect 23224 32678 23230 32734
rect 23951 32585 24064 32591
rect 23103 32472 23951 32585
rect 23103 32437 23216 32472
rect 23951 32466 24064 32472
rect 23097 32425 23221 32437
rect 23444 32430 23500 32436
rect 23097 32313 23103 32425
rect 23215 32313 23221 32425
rect 23346 32374 23352 32430
rect 23408 32374 23414 32430
rect 23444 32368 23500 32374
rect 23097 32301 23221 32313
rect 23846 32308 23852 32364
rect 23908 32358 24790 32364
rect 23908 32314 24734 32358
rect 24778 32314 24790 32358
rect 23908 32308 24790 32314
rect 23254 32130 23260 32187
rect 23316 32130 23322 32187
rect 23444 32112 23500 32168
rect 23159 31947 23221 31959
rect 20659 31941 23165 31947
rect 20659 31903 20671 31941
rect 20709 31903 23165 31941
rect 20659 31897 23165 31903
rect 23215 31897 23221 31947
rect 23159 31891 23221 31897
rect 23159 31885 23215 31891
rect 23346 31889 23352 31945
rect 23408 31889 23414 31945
rect 23165 31863 23215 31885
rect 23530 31868 23536 31924
rect 23592 31868 23598 31924
rect 23945 31876 23951 31989
rect 24064 31945 24070 31989
rect 24068 31936 24074 31945
rect 26045 31936 26103 31942
rect 24068 31902 26057 31936
rect 26091 31902 26103 31936
rect 24068 31893 24074 31902
rect 26045 31896 26103 31902
rect 24064 31876 24070 31893
rect 23173 31800 23214 31863
rect 23863 31806 23915 31812
rect 23173 31759 23863 31800
rect 23863 31748 23915 31754
rect 23162 31588 23168 31644
rect 23224 31588 23230 31644
rect 22511 29582 23352 29583
rect 22511 29527 22616 29582
rect 22610 29526 22616 29527
rect 22672 29527 23352 29582
rect 23408 29527 23415 29583
rect 22672 29526 22678 29527
rect 23162 29414 23168 29470
rect 23224 29414 23230 29470
rect 23951 29321 24064 29327
rect 23103 29208 23951 29321
rect 23103 29173 23216 29208
rect 23951 29202 24064 29208
rect 23097 29161 23221 29173
rect 23444 29166 23500 29172
rect 23097 29049 23103 29161
rect 23215 29049 23221 29161
rect 23346 29110 23352 29166
rect 23408 29110 23414 29166
rect 23444 29104 23500 29110
rect 23097 29037 23221 29049
rect 23846 29044 23852 29100
rect 23908 29094 24790 29100
rect 23908 29050 24734 29094
rect 24778 29050 24790 29094
rect 23908 29044 24790 29050
rect 23254 28866 23260 28923
rect 23316 28866 23322 28923
rect 23444 28848 23500 28904
rect 23159 28683 23221 28695
rect 20659 28677 23165 28683
rect 20659 28639 20671 28677
rect 20709 28639 23165 28677
rect 20659 28633 23165 28639
rect 23215 28633 23221 28683
rect 23159 28627 23221 28633
rect 23159 28621 23215 28627
rect 23346 28625 23352 28681
rect 23408 28625 23414 28681
rect 23165 28599 23215 28621
rect 23530 28604 23536 28660
rect 23592 28604 23598 28660
rect 23945 28612 23951 28725
rect 24064 28681 24070 28725
rect 24068 28672 24074 28681
rect 26045 28672 26103 28678
rect 24068 28638 26057 28672
rect 26091 28638 26103 28672
rect 24068 28629 24074 28638
rect 26045 28632 26103 28638
rect 24064 28612 24070 28629
rect 23173 28536 23214 28599
rect 23863 28542 23915 28548
rect 23173 28495 23863 28536
rect 23863 28484 23915 28490
rect 23162 28324 23168 28380
rect 23224 28324 23230 28380
rect 22511 26318 23352 26319
rect 22511 26263 22708 26318
rect 22702 26262 22708 26263
rect 22764 26263 23352 26318
rect 23408 26263 23415 26319
rect 22764 26262 22770 26263
rect 23162 26150 23168 26206
rect 23224 26150 23230 26206
rect 23951 26057 24064 26063
rect 23103 25944 23951 26057
rect 23103 25909 23216 25944
rect 23951 25938 24064 25944
rect 23097 25897 23221 25909
rect 23444 25902 23500 25908
rect 23097 25785 23103 25897
rect 23215 25785 23221 25897
rect 23346 25846 23352 25902
rect 23408 25846 23414 25902
rect 23444 25840 23500 25846
rect 23097 25773 23221 25785
rect 23846 25780 23852 25836
rect 23908 25830 24790 25836
rect 23908 25786 24734 25830
rect 24778 25786 24790 25830
rect 23908 25780 24790 25786
rect 23254 25602 23260 25659
rect 23316 25602 23322 25659
rect 23444 25584 23500 25640
rect 23159 25419 23221 25431
rect 20659 25413 23165 25419
rect 20659 25375 20671 25413
rect 20709 25375 23165 25413
rect 20659 25369 23165 25375
rect 23215 25369 23221 25419
rect 23159 25363 23221 25369
rect 23159 25357 23215 25363
rect 23346 25361 23352 25417
rect 23408 25361 23414 25417
rect 23165 25335 23215 25357
rect 23530 25340 23536 25396
rect 23592 25340 23598 25396
rect 23945 25348 23951 25461
rect 24064 25417 24070 25461
rect 24068 25408 24074 25417
rect 26045 25408 26103 25414
rect 24068 25374 26057 25408
rect 26091 25374 26103 25408
rect 24068 25365 24074 25374
rect 26045 25368 26103 25374
rect 24064 25348 24070 25365
rect 23173 25272 23214 25335
rect 23863 25278 23915 25284
rect 23173 25231 23863 25272
rect 23863 25220 23915 25226
rect 23162 25060 23168 25116
rect 23224 25060 23230 25116
rect 1763 23243 1815 23249
rect 438 23184 444 23243
rect 503 23209 1769 23243
rect 1803 23209 1815 23243
rect 503 23184 509 23209
rect 1763 23203 1815 23209
rect 22511 23054 23352 23055
rect 22511 22999 22800 23054
rect 22794 22998 22800 22999
rect 22856 22999 23352 23054
rect 23408 22999 23415 23055
rect 22856 22998 22862 22999
rect 23162 22886 23168 22942
rect 23224 22886 23230 22942
rect 23951 22793 24064 22799
rect 23103 22680 23951 22793
rect 23103 22645 23216 22680
rect 23951 22674 24064 22680
rect 23097 22633 23221 22645
rect 23444 22638 23500 22644
rect 23097 22521 23103 22633
rect 23215 22521 23221 22633
rect 23346 22582 23352 22638
rect 23408 22582 23414 22638
rect 23444 22576 23500 22582
rect 23097 22509 23221 22521
rect 23846 22516 23852 22572
rect 23908 22566 24790 22572
rect 23908 22522 24734 22566
rect 24778 22522 24790 22566
rect 23908 22516 24790 22522
rect 23254 22338 23260 22395
rect 23316 22338 23322 22395
rect 23444 22320 23500 22376
rect 23159 22155 23221 22167
rect 20659 22149 23165 22155
rect 20659 22111 20671 22149
rect 20709 22111 23165 22149
rect 20659 22105 23165 22111
rect 23215 22105 23221 22155
rect 23159 22099 23221 22105
rect 23159 22093 23215 22099
rect 23346 22097 23352 22153
rect 23408 22097 23414 22153
rect 23165 22071 23215 22093
rect 23530 22076 23536 22132
rect 23592 22076 23598 22132
rect 23945 22084 23951 22197
rect 24064 22153 24070 22197
rect 24068 22144 24074 22153
rect 26045 22144 26103 22150
rect 24068 22110 26057 22144
rect 26091 22110 26103 22144
rect 24068 22101 24074 22110
rect 26045 22104 26103 22110
rect 24064 22084 24070 22101
rect 23173 22008 23214 22071
rect 23863 22014 23915 22020
rect 23173 21967 23863 22008
rect 23863 21956 23915 21962
rect 23162 21796 23168 21852
rect 23224 21796 23230 21852
rect 436 20413 510 20419
rect 430 20351 436 20413
rect 510 20351 516 20413
rect 430 20345 442 20351
rect 504 20345 516 20351
rect 430 20339 516 20345
rect 1763 19979 1815 19985
rect 438 19920 444 19979
rect 503 19945 1769 19979
rect 1803 19945 1815 19979
rect 503 19920 509 19945
rect 1763 19939 1815 19945
rect 22511 19790 23352 19791
rect 22511 19735 22892 19790
rect 22886 19734 22892 19735
rect 22948 19735 23352 19790
rect 23408 19735 23415 19791
rect 22948 19734 22954 19735
rect 23162 19622 23168 19678
rect 23224 19622 23230 19678
rect 23951 19529 24064 19535
rect 23103 19416 23951 19529
rect 23103 19381 23216 19416
rect 23951 19410 24064 19416
rect 23097 19369 23221 19381
rect 23444 19374 23500 19380
rect 23097 19257 23103 19369
rect 23215 19257 23221 19369
rect 23346 19318 23352 19374
rect 23408 19318 23414 19374
rect 23444 19312 23500 19318
rect 23097 19245 23221 19257
rect 23846 19252 23852 19308
rect 23908 19302 24790 19308
rect 23908 19258 24734 19302
rect 24778 19258 24790 19302
rect 23908 19252 24790 19258
rect 23254 19074 23260 19131
rect 23316 19074 23322 19131
rect 23444 19056 23500 19112
rect 23159 18891 23221 18903
rect 20659 18885 23165 18891
rect 20659 18847 20671 18885
rect 20709 18847 23165 18885
rect 20659 18841 23165 18847
rect 23215 18841 23221 18891
rect 23159 18835 23221 18841
rect 23159 18829 23215 18835
rect 23346 18833 23352 18889
rect 23408 18833 23414 18889
rect 23165 18807 23215 18829
rect 23530 18812 23536 18868
rect 23592 18812 23598 18868
rect 23945 18820 23951 18933
rect 24064 18889 24070 18933
rect 24068 18880 24074 18889
rect 26045 18880 26103 18886
rect 24068 18846 26057 18880
rect 26091 18846 26103 18880
rect 24068 18837 24074 18846
rect 26045 18840 26103 18846
rect 24064 18820 24070 18837
rect 23173 18744 23214 18807
rect 23863 18750 23915 18756
rect 23173 18703 23863 18744
rect 23863 18692 23915 18698
rect 23162 18532 23168 18588
rect 23224 18532 23230 18588
rect 436 17149 510 17155
rect 430 17087 436 17149
rect 510 17087 516 17149
rect 430 17081 442 17087
rect 504 17081 516 17087
rect 430 17075 516 17081
rect 1763 16715 1815 16721
rect 438 16656 444 16715
rect 503 16681 1769 16715
rect 1803 16681 1815 16715
rect 503 16656 509 16681
rect 1763 16675 1815 16681
rect 22978 16527 22984 16528
rect 22511 16472 22984 16527
rect 23040 16527 23046 16528
rect 23040 16472 23352 16527
rect 22511 16471 23352 16472
rect 23408 16471 23415 16527
rect 23162 16358 23168 16414
rect 23224 16358 23230 16414
rect 23951 16265 24064 16271
rect 23103 16152 23951 16265
rect 23103 16117 23216 16152
rect 23951 16146 24064 16152
rect 23097 16105 23221 16117
rect 23444 16110 23500 16116
rect 23097 15993 23103 16105
rect 23215 15993 23221 16105
rect 23346 16054 23352 16110
rect 23408 16054 23414 16110
rect 23444 16048 23500 16054
rect 23097 15981 23221 15993
rect 23846 15988 23852 16044
rect 23908 16038 24790 16044
rect 23908 15994 24734 16038
rect 24778 15994 24790 16038
rect 23908 15988 24790 15994
rect 23254 15810 23260 15867
rect 23316 15810 23322 15867
rect 23444 15792 23500 15848
rect 23159 15627 23221 15639
rect 20659 15621 23165 15627
rect 20659 15583 20671 15621
rect 20709 15583 23165 15621
rect 20659 15577 23165 15583
rect 23215 15577 23221 15627
rect 23159 15571 23221 15577
rect 23159 15565 23215 15571
rect 23346 15569 23352 15625
rect 23408 15569 23414 15625
rect 23165 15543 23215 15565
rect 23530 15548 23536 15604
rect 23592 15548 23598 15604
rect 23945 15556 23951 15669
rect 24064 15625 24070 15669
rect 24068 15616 24074 15625
rect 26045 15616 26103 15622
rect 24068 15582 26057 15616
rect 26091 15582 26103 15616
rect 24068 15573 24074 15582
rect 26045 15576 26103 15582
rect 24064 15556 24070 15573
rect 23173 15480 23214 15543
rect 23863 15486 23915 15492
rect 23173 15439 23863 15480
rect 23863 15428 23915 15434
rect 23162 15268 23168 15324
rect 23224 15268 23230 15324
rect 436 13885 510 13891
rect 430 13823 436 13885
rect 510 13823 516 13885
rect 430 13817 442 13823
rect 504 13817 516 13823
rect 430 13811 516 13817
rect 1763 13451 1815 13457
rect 438 13392 444 13451
rect 503 13417 1769 13451
rect 1803 13417 1815 13451
rect 503 13392 509 13417
rect 1763 13411 1815 13417
rect 22511 13260 23352 13263
rect 22511 13207 23076 13260
rect 23070 13204 23076 13207
rect 23132 13207 23352 13260
rect 23408 13207 23415 13263
rect 23132 13204 23138 13207
rect 23162 13094 23168 13150
rect 23224 13094 23230 13150
rect 23951 13001 24064 13007
rect 23103 12888 23951 13001
rect 23103 12853 23216 12888
rect 23951 12882 24064 12888
rect 23097 12841 23221 12853
rect 23444 12846 23500 12852
rect 23097 12729 23103 12841
rect 23215 12729 23221 12841
rect 23346 12790 23352 12846
rect 23408 12790 23414 12846
rect 23444 12784 23500 12790
rect 23097 12717 23221 12729
rect 23846 12724 23852 12780
rect 23908 12774 24790 12780
rect 23908 12730 24734 12774
rect 24778 12730 24790 12774
rect 23908 12724 24790 12730
rect 23254 12547 23260 12603
rect 23316 12547 23322 12603
rect 23444 12528 23500 12584
rect 11884 12008 11890 12064
rect 11946 12008 11952 12064
rect 11099 11824 11105 11884
rect 11165 11824 11171 11884
rect 10620 11811 10706 11823
rect 10620 11805 10626 11811
rect 10700 11805 10706 11811
rect 9981 11746 10067 11752
rect 6024 11617 6030 11724
rect 6137 11703 9894 11724
rect 6137 11637 9807 11703
rect 9873 11637 9894 11703
rect 9981 11678 9993 11746
rect 10061 11740 10246 11746
rect 10061 11684 10178 11740
rect 10234 11684 10246 11740
rect 12667 11808 12741 11814
rect 11400 11798 11473 11804
rect 11400 11795 11412 11798
rect 11461 11795 11473 11798
rect 11400 11743 11406 11795
rect 11467 11743 11473 11795
rect 11523 11760 11575 11766
rect 11406 11737 11467 11743
rect 10620 11725 10706 11731
rect 11651 11731 11657 11801
rect 11727 11731 11733 11801
rect 12667 11752 12679 11808
rect 12735 11752 23444 11808
rect 23500 11752 23729 11808
rect 12447 11746 12516 11752
rect 12667 11746 12741 11752
rect 11523 11702 11575 11708
rect 12447 11701 12459 11746
rect 12504 11701 12516 11746
rect 12447 11695 12516 11701
rect 10061 11678 10246 11684
rect 9981 11677 10067 11678
rect 9987 11672 10067 11677
rect 6137 11617 9894 11637
rect 12459 11667 12504 11695
rect 23528 11670 23534 11674
rect 12544 11667 23534 11670
rect 12459 11625 23534 11667
rect 23528 11622 23534 11625
rect 23586 11670 23592 11674
rect 23586 11625 23729 11670
rect 23586 11622 23592 11625
rect 12051 11461 12057 11517
rect 12113 11461 12119 11517
rect 11890 11126 11946 11132
rect 11946 11070 23168 11126
rect 23224 11070 23230 11126
rect 11890 11064 11946 11070
rect 12051 10959 12057 11015
rect 12113 10959 23260 11015
rect 23316 10959 23322 11015
rect 436 10621 510 10627
rect 430 10559 436 10621
rect 510 10559 516 10621
rect 430 10553 442 10559
rect 504 10553 516 10559
rect 430 10547 516 10553
rect 1763 10187 1815 10193
rect 438 10128 444 10187
rect 503 10153 1769 10187
rect 1803 10153 1815 10187
rect 503 10128 509 10153
rect 1763 10147 1815 10153
rect 19794 10053 19852 10059
rect 19852 9995 26888 10053
rect 26946 9995 26952 10053
rect 19794 9989 19852 9995
rect 19516 9866 19522 9924
rect 19580 9866 27164 9924
rect 27222 9866 27228 9924
rect 19247 9775 19305 9781
rect 19305 9717 27439 9775
rect 27497 9717 27503 9775
rect 19247 9711 19305 9717
rect 18956 9545 18962 9603
rect 19020 9545 27714 9603
rect 27772 9545 27778 9603
rect 18417 9377 18423 9435
rect 18481 9377 28271 9435
rect 28329 9377 28335 9435
rect 18297 9277 18303 9335
rect 18361 9277 28391 9335
rect 28449 9277 28455 9335
rect 18174 9150 18180 9208
rect 18238 9150 28511 9208
rect 28569 9150 28575 9208
rect 18055 9037 18061 9095
rect 18119 9037 28631 9095
rect 28689 9037 28695 9095
rect 436 7357 510 7363
rect 430 7295 436 7357
rect 510 7295 516 7357
rect 430 7289 442 7295
rect 504 7289 516 7295
rect 430 7283 516 7289
rect 1763 6923 1815 6929
rect 438 6864 444 6923
rect 503 6889 1769 6923
rect 1803 6889 1815 6923
rect 503 6864 509 6889
rect 1763 6883 1815 6889
rect 436 4093 510 4099
rect 430 4031 436 4093
rect 510 4031 516 4093
rect 430 4025 442 4031
rect 504 4025 516 4031
rect 430 4019 516 4025
rect 1763 3659 1815 3665
rect 438 3600 444 3659
rect 503 3625 1769 3659
rect 1803 3625 1815 3659
rect 503 3600 509 3625
rect 1763 3619 1815 3625
rect 436 829 510 835
rect 430 767 436 829
rect 510 767 516 829
rect 430 761 442 767
rect 504 761 516 767
rect 430 755 516 761
rect 11523 369 11575 375
rect 10725 317 10731 369
rect 10783 359 10789 369
rect 10783 327 11523 359
rect 10783 317 10789 327
rect 11523 311 11575 317
rect 10803 231 10809 283
rect 10861 281 10867 283
rect 11405 281 11411 282
rect 10861 232 11411 281
rect 10861 231 10867 232
rect 11405 230 11411 232
rect 11463 230 11469 282
rect -424 16 78 112
rect 8949 108 8980 112
<< via1 >>
rect 23260 35394 23316 35450
rect 23352 35203 23408 35209
rect 23352 35159 23358 35203
rect 23358 35159 23402 35203
rect 23402 35159 23408 35203
rect 23352 35153 23408 35159
rect 23536 35182 23592 35188
rect 23536 35138 23542 35182
rect 23542 35138 23586 35182
rect 23586 35138 23592 35182
rect 23536 35132 23592 35138
rect 23951 35209 24064 35253
rect 23951 35157 24068 35209
rect 23951 35140 24064 35157
rect 23863 35018 23915 35070
rect 23168 34852 23224 34908
rect 22524 32792 22580 32848
rect 23352 32791 23408 32847
rect 23168 32678 23224 32734
rect 23951 32472 24064 32585
rect 23352 32424 23408 32430
rect 23352 32380 23358 32424
rect 23358 32380 23402 32424
rect 23402 32380 23408 32424
rect 23352 32374 23408 32380
rect 23444 32424 23500 32430
rect 23444 32380 23450 32424
rect 23450 32380 23494 32424
rect 23494 32380 23500 32424
rect 23444 32374 23500 32380
rect 23852 32308 23908 32364
rect 23260 32130 23316 32187
rect 23352 31939 23408 31945
rect 23352 31895 23358 31939
rect 23358 31895 23402 31939
rect 23402 31895 23408 31939
rect 23352 31889 23408 31895
rect 23536 31918 23592 31924
rect 23536 31874 23542 31918
rect 23542 31874 23586 31918
rect 23586 31874 23592 31918
rect 23536 31868 23592 31874
rect 23951 31945 24064 31989
rect 23951 31893 24068 31945
rect 23951 31876 24064 31893
rect 23863 31754 23915 31806
rect 23168 31588 23224 31644
rect 22616 29526 22672 29582
rect 23352 29527 23408 29583
rect 23168 29414 23224 29470
rect 23951 29208 24064 29321
rect 23352 29160 23408 29166
rect 23352 29116 23358 29160
rect 23358 29116 23402 29160
rect 23402 29116 23408 29160
rect 23352 29110 23408 29116
rect 23444 29160 23500 29166
rect 23444 29116 23450 29160
rect 23450 29116 23494 29160
rect 23494 29116 23500 29160
rect 23444 29110 23500 29116
rect 23852 29044 23908 29100
rect 23260 28866 23316 28923
rect 23352 28675 23408 28681
rect 23352 28631 23358 28675
rect 23358 28631 23402 28675
rect 23402 28631 23408 28675
rect 23352 28625 23408 28631
rect 23536 28654 23592 28660
rect 23536 28610 23542 28654
rect 23542 28610 23586 28654
rect 23586 28610 23592 28654
rect 23536 28604 23592 28610
rect 23951 28681 24064 28725
rect 23951 28629 24068 28681
rect 23951 28612 24064 28629
rect 23863 28490 23915 28542
rect 23168 28324 23224 28380
rect 22708 26262 22764 26318
rect 23352 26263 23408 26319
rect 23168 26150 23224 26206
rect 23951 25944 24064 26057
rect 23352 25896 23408 25902
rect 23352 25852 23358 25896
rect 23358 25852 23402 25896
rect 23402 25852 23408 25896
rect 23352 25846 23408 25852
rect 23444 25896 23500 25902
rect 23444 25852 23450 25896
rect 23450 25852 23494 25896
rect 23494 25852 23500 25896
rect 23444 25846 23500 25852
rect 23852 25780 23908 25836
rect 23260 25602 23316 25659
rect 23352 25411 23408 25417
rect 23352 25367 23358 25411
rect 23358 25367 23402 25411
rect 23402 25367 23408 25411
rect 23352 25361 23408 25367
rect 23536 25390 23592 25396
rect 23536 25346 23542 25390
rect 23542 25346 23586 25390
rect 23586 25346 23592 25390
rect 23536 25340 23592 25346
rect 23951 25417 24064 25461
rect 23951 25365 24068 25417
rect 23951 25348 24064 25365
rect 23863 25226 23915 25278
rect 23168 25060 23224 25116
rect 444 23184 503 23243
rect 22800 22998 22856 23054
rect 23352 22999 23408 23055
rect 23168 22886 23224 22942
rect 23951 22680 24064 22793
rect 23352 22632 23408 22638
rect 23352 22588 23358 22632
rect 23358 22588 23402 22632
rect 23402 22588 23408 22632
rect 23352 22582 23408 22588
rect 23444 22632 23500 22638
rect 23444 22588 23450 22632
rect 23450 22588 23494 22632
rect 23494 22588 23500 22632
rect 23444 22582 23500 22588
rect 23852 22516 23908 22572
rect 23260 22338 23316 22395
rect 23352 22147 23408 22153
rect 23352 22103 23358 22147
rect 23358 22103 23402 22147
rect 23402 22103 23408 22147
rect 23352 22097 23408 22103
rect 23536 22126 23592 22132
rect 23536 22082 23542 22126
rect 23542 22082 23586 22126
rect 23586 22082 23592 22126
rect 23536 22076 23592 22082
rect 23951 22153 24064 22197
rect 23951 22101 24068 22153
rect 23951 22084 24064 22101
rect 23863 21962 23915 22014
rect 23168 21796 23224 21852
rect 436 20407 510 20413
rect 436 20351 442 20407
rect 442 20351 504 20407
rect 504 20351 510 20407
rect 444 19920 503 19979
rect 22892 19734 22948 19790
rect 23352 19735 23408 19791
rect 23168 19622 23224 19678
rect 23951 19416 24064 19529
rect 23352 19368 23408 19374
rect 23352 19324 23358 19368
rect 23358 19324 23402 19368
rect 23402 19324 23408 19368
rect 23352 19318 23408 19324
rect 23444 19368 23500 19374
rect 23444 19324 23450 19368
rect 23450 19324 23494 19368
rect 23494 19324 23500 19368
rect 23444 19318 23500 19324
rect 23852 19252 23908 19308
rect 23260 19074 23316 19131
rect 23352 18883 23408 18889
rect 23352 18839 23358 18883
rect 23358 18839 23402 18883
rect 23402 18839 23408 18883
rect 23352 18833 23408 18839
rect 23536 18862 23592 18868
rect 23536 18818 23542 18862
rect 23542 18818 23586 18862
rect 23586 18818 23592 18862
rect 23536 18812 23592 18818
rect 23951 18889 24064 18933
rect 23951 18837 24068 18889
rect 23951 18820 24064 18837
rect 23863 18698 23915 18750
rect 23168 18532 23224 18588
rect 436 17143 510 17149
rect 436 17087 442 17143
rect 442 17087 504 17143
rect 504 17087 510 17143
rect 444 16656 503 16715
rect 22984 16472 23040 16528
rect 23352 16471 23408 16527
rect 23168 16358 23224 16414
rect 23951 16152 24064 16265
rect 23352 16104 23408 16110
rect 23352 16060 23358 16104
rect 23358 16060 23402 16104
rect 23402 16060 23408 16104
rect 23352 16054 23408 16060
rect 23444 16104 23500 16110
rect 23444 16060 23450 16104
rect 23450 16060 23494 16104
rect 23494 16060 23500 16104
rect 23444 16054 23500 16060
rect 23852 15988 23908 16044
rect 23260 15810 23316 15867
rect 23352 15619 23408 15625
rect 23352 15575 23358 15619
rect 23358 15575 23402 15619
rect 23402 15575 23408 15619
rect 23352 15569 23408 15575
rect 23536 15598 23592 15604
rect 23536 15554 23542 15598
rect 23542 15554 23586 15598
rect 23586 15554 23592 15598
rect 23536 15548 23592 15554
rect 23951 15625 24064 15669
rect 23951 15573 24068 15625
rect 23951 15556 24064 15573
rect 23863 15434 23915 15486
rect 23168 15268 23224 15324
rect 436 13879 510 13885
rect 436 13823 442 13879
rect 442 13823 504 13879
rect 504 13823 510 13879
rect 444 13392 503 13451
rect 23076 13204 23132 13260
rect 23352 13207 23408 13263
rect 23168 13094 23224 13150
rect 23951 12888 24064 13001
rect 23352 12840 23408 12846
rect 23352 12796 23358 12840
rect 23358 12796 23402 12840
rect 23402 12796 23408 12840
rect 23352 12790 23408 12796
rect 23444 12840 23500 12846
rect 23444 12796 23450 12840
rect 23450 12796 23494 12840
rect 23494 12796 23500 12840
rect 23444 12790 23500 12796
rect 23852 12724 23908 12780
rect 23260 12547 23316 12603
rect 11890 12008 11946 12064
rect 11105 11878 11165 11884
rect 11105 11830 11111 11878
rect 11111 11830 11159 11878
rect 11159 11830 11165 11878
rect 11105 11824 11165 11830
rect 6030 11617 6137 11724
rect 10620 11737 10626 11805
rect 10626 11737 10700 11805
rect 10700 11737 10706 11805
rect 11406 11749 11412 11795
rect 11412 11749 11461 11795
rect 11461 11749 11467 11795
rect 11406 11743 11467 11749
rect 11523 11751 11575 11760
rect 10620 11731 10706 11737
rect 11523 11717 11532 11751
rect 11532 11717 11566 11751
rect 11566 11717 11575 11751
rect 11657 11795 11727 11801
rect 11657 11737 11663 11795
rect 11663 11737 11721 11795
rect 11721 11737 11727 11795
rect 11657 11731 11727 11737
rect 23444 11752 23500 11808
rect 11523 11708 11575 11717
rect 23534 11622 23586 11674
rect 12057 11461 12113 11517
rect 11890 11070 11946 11126
rect 23168 11070 23224 11126
rect 12057 10959 12113 11015
rect 23260 10959 23316 11015
rect 436 10615 510 10621
rect 436 10559 442 10615
rect 442 10559 504 10615
rect 504 10559 510 10615
rect 444 10128 503 10187
rect 19794 9995 19852 10053
rect 26888 9995 26946 10053
rect 19522 9866 19580 9924
rect 27164 9866 27222 9924
rect 19247 9717 19305 9775
rect 27439 9717 27497 9775
rect 18962 9545 19020 9603
rect 27714 9545 27772 9603
rect 18423 9377 18481 9435
rect 28271 9377 28329 9435
rect 18303 9277 18361 9335
rect 28391 9277 28449 9335
rect 18180 9150 18238 9208
rect 28511 9150 28569 9208
rect 18061 9037 18119 9095
rect 28631 9037 28689 9095
rect 436 7351 510 7357
rect 436 7295 442 7351
rect 442 7295 504 7351
rect 504 7295 510 7351
rect 444 6864 503 6923
rect 436 4087 510 4093
rect 436 4031 442 4087
rect 442 4031 504 4087
rect 504 4031 510 4087
rect 444 3600 503 3659
rect 436 823 510 829
rect 436 767 442 823
rect 442 767 504 823
rect 504 767 510 823
rect 10731 317 10783 369
rect 11523 317 11575 369
rect 10809 231 10861 283
rect 11411 230 11463 282
<< metal2 >>
rect 16333 34122 16422 35472
rect 23168 34908 23224 35472
rect 22524 32848 22580 32855
rect 444 23243 503 23249
rect 444 20413 503 23184
rect 6046 22576 6142 23504
rect -276 20351 436 20413
rect 510 20351 516 20413
rect -276 16 -217 20351
rect 444 20339 503 20351
rect 444 19979 503 19985
rect 444 17149 503 19920
rect -156 17087 436 17149
rect 510 17087 516 17149
rect -156 16 -97 17087
rect 444 17075 503 17087
rect 444 16715 503 16721
rect 444 13885 503 16656
rect -36 13823 436 13885
rect 510 13823 516 13885
rect -36 16 23 13823
rect 444 13811 503 13823
rect 444 13451 503 13457
rect 444 10621 503 13392
rect 11890 12064 11946 12070
rect 11105 11884 11165 11890
rect 10614 11731 10620 11805
rect 10706 11731 10712 11805
rect 6030 11724 6137 11730
rect 6030 11611 6137 11617
rect 84 10559 436 10621
rect 510 10559 516 10621
rect 84 16 143 10559
rect 444 10547 503 10559
rect 444 10187 503 10193
rect 444 7357 503 10128
rect 204 7295 436 7357
rect 510 7295 516 7357
rect 204 16 263 7295
rect 444 7283 503 7295
rect 444 6923 503 6929
rect 444 4093 503 6864
rect 324 4031 436 4093
rect 510 4031 516 4093
rect 324 16 383 4031
rect 444 4019 503 4031
rect 444 3659 503 3665
rect 444 829 503 3600
rect 430 767 436 829
rect 510 767 516 829
rect 444 16 503 767
rect 2600 16 2658 112
rect 2876 16 2934 112
rect 3151 16 3209 112
rect 3426 16 3484 112
rect 3983 16 4041 112
rect 4103 16 4161 112
rect 4223 16 4281 112
rect 4343 16 4401 112
rect 10626 16 10700 11731
rect 10731 369 10783 375
rect 10731 311 10783 317
rect 10741 16 10773 311
rect 10809 283 10861 289
rect 10809 225 10861 231
rect 10811 16 10860 225
rect 11105 16 11165 11824
rect 11657 11801 11727 11807
rect 11400 11743 11406 11795
rect 11467 11743 11473 11795
rect 11412 288 11461 11743
rect 11517 11708 11523 11760
rect 11575 11708 11581 11760
rect 11657 11725 11727 11731
rect 11533 369 11565 11708
rect 11517 317 11523 369
rect 11575 317 11581 369
rect 11411 282 11463 288
rect 11411 224 11463 230
rect 11663 16 11723 11725
rect 11890 11126 11946 12008
rect 12057 11517 12113 11523
rect 11884 11070 11890 11126
rect 11946 11070 11952 11126
rect 11890 16 11946 11070
rect 12057 11015 12113 11461
rect 12057 16 12113 10959
rect 18067 9101 18125 12180
rect 18187 9214 18245 12101
rect 18307 9341 18365 12081
rect 18427 9441 18485 12142
rect 18984 9609 19042 12073
rect 19259 9775 19317 12176
rect 19534 9930 19592 12065
rect 19810 10053 19868 12103
rect 19788 9995 19794 10053
rect 19852 9995 19868 10053
rect 19522 9924 19592 9930
rect 19580 9866 19592 9924
rect 19522 9860 19592 9866
rect 19241 9717 19247 9775
rect 19305 9717 19317 9775
rect 18962 9603 19042 9609
rect 19020 9545 19042 9603
rect 18962 9539 19042 9545
rect 18423 9435 18485 9441
rect 18481 9377 18485 9435
rect 18423 9371 18485 9377
rect 18303 9335 18365 9341
rect 18361 9277 18365 9335
rect 18303 9271 18365 9277
rect 18180 9208 18245 9214
rect 18238 9150 18245 9208
rect 18180 9144 18245 9150
rect 18061 9095 18125 9101
rect 18119 9037 18125 9095
rect 18061 9031 18125 9037
rect 18067 16 18125 9031
rect 18187 16 18245 9144
rect 18307 16 18365 9271
rect 18427 16 18485 9371
rect 18984 16 19042 9539
rect 19259 16 19317 9717
rect 19534 16 19592 9860
rect 19810 16 19868 9995
rect 22524 16 22580 32792
rect 23168 32734 23224 34852
rect 23168 31644 23224 32678
rect 22616 29582 22672 29590
rect 22616 16 22672 29526
rect 23168 29470 23224 31588
rect 23168 28380 23224 29414
rect 22708 26318 22764 26325
rect 22708 16 22764 26262
rect 23168 26206 23224 28324
rect 23168 25116 23224 26150
rect 22800 23054 22856 23061
rect 22800 16 22856 22998
rect 23168 22942 23224 25060
rect 23168 21852 23224 22886
rect 22892 19790 22948 19798
rect 22892 16 22948 19734
rect 23168 19678 23224 21796
rect 23168 18588 23224 19622
rect 22984 16528 23040 16537
rect 22984 16 23040 16472
rect 23168 16414 23224 18532
rect 23168 15324 23224 16358
rect 23076 13260 23132 13266
rect 23076 16 23132 13204
rect 23168 13150 23224 15268
rect 23168 11126 23224 13094
rect 23168 11064 23224 11070
rect 23260 35450 23316 35472
rect 23260 32187 23316 35394
rect 23352 35209 23408 35215
rect 23352 32847 23408 35153
rect 23352 32430 23408 32791
rect 23444 32430 23500 35376
rect 23536 35188 23592 35376
rect 23438 32374 23444 32430
rect 23500 32374 23506 32430
rect 23352 32368 23408 32374
rect 23260 28923 23316 32130
rect 23352 31945 23408 31951
rect 23352 29583 23408 31889
rect 23352 29166 23408 29527
rect 23444 29166 23500 32374
rect 23536 31924 23592 35132
rect 23951 35253 24064 35259
rect 24064 35209 24068 35215
rect 24064 35151 24068 35157
rect 23852 35070 23908 35076
rect 23852 35018 23863 35070
rect 23915 35018 23921 35070
rect 23852 32364 23908 35018
rect 23951 32585 24064 35140
rect 30334 34175 30423 35472
rect 23945 32472 23951 32585
rect 24064 32472 24070 32585
rect 23852 32302 23908 32308
rect 23438 29110 23444 29166
rect 23500 29110 23506 29166
rect 23352 29104 23408 29110
rect 23260 25659 23316 28866
rect 23352 28681 23408 28687
rect 23352 26319 23408 28625
rect 23352 25902 23408 26263
rect 23444 25902 23500 29110
rect 23536 28660 23592 31868
rect 23951 31989 24064 31995
rect 24064 31945 24068 31951
rect 24064 31887 24068 31893
rect 23852 31806 23908 31812
rect 23852 31754 23863 31806
rect 23915 31754 23921 31806
rect 23852 29100 23908 31754
rect 23951 29321 24064 31876
rect 23945 29208 23951 29321
rect 24064 29208 24070 29321
rect 23852 29038 23908 29044
rect 23438 25846 23444 25902
rect 23500 25846 23506 25902
rect 23352 25840 23408 25846
rect 23260 22395 23316 25602
rect 23352 25417 23408 25423
rect 23352 23055 23408 25361
rect 23352 22638 23408 22999
rect 23444 22638 23500 25846
rect 23536 25396 23592 28604
rect 23951 28725 24064 28731
rect 24064 28681 24068 28687
rect 24064 28623 24068 28629
rect 23852 28542 23908 28548
rect 23852 28490 23863 28542
rect 23915 28490 23921 28542
rect 23852 25836 23908 28490
rect 23951 26057 24064 28612
rect 23945 25944 23951 26057
rect 24064 25944 24070 26057
rect 23852 25774 23908 25780
rect 23438 22582 23444 22638
rect 23500 22582 23506 22638
rect 23352 22576 23408 22582
rect 23260 19131 23316 22338
rect 23352 22153 23408 22159
rect 23352 19791 23408 22097
rect 23352 19374 23408 19735
rect 23444 19374 23500 22582
rect 23536 22132 23592 25340
rect 23951 25461 24064 25467
rect 24064 25417 24068 25423
rect 24064 25359 24068 25365
rect 23852 25278 23908 25284
rect 23852 25226 23863 25278
rect 23915 25226 23921 25278
rect 23852 22572 23908 25226
rect 23951 22793 24064 25348
rect 23945 22680 23951 22793
rect 24064 22680 24070 22793
rect 23852 22510 23908 22516
rect 23438 19318 23444 19374
rect 23500 19318 23506 19374
rect 23352 19312 23408 19318
rect 23260 15867 23316 19074
rect 23352 18889 23408 18895
rect 23352 16527 23408 18833
rect 23352 16110 23408 16471
rect 23444 16110 23500 19318
rect 23536 18868 23592 22076
rect 23951 22197 24064 22203
rect 24064 22153 24068 22159
rect 24064 22095 24068 22101
rect 23852 22014 23908 22020
rect 23852 21962 23863 22014
rect 23915 21962 23921 22014
rect 23852 19308 23908 21962
rect 23951 19529 24064 22084
rect 23945 19416 23951 19529
rect 24064 19416 24070 19529
rect 23852 19246 23908 19252
rect 23438 16054 23444 16110
rect 23500 16054 23506 16110
rect 23352 16048 23408 16054
rect 23260 12603 23316 15810
rect 23352 15625 23408 15631
rect 23352 13263 23408 15569
rect 23352 12846 23408 13207
rect 23444 12846 23500 16054
rect 23536 15604 23592 18812
rect 23951 18933 24064 18939
rect 24064 18889 24068 18895
rect 24064 18831 24068 18837
rect 23852 18750 23908 18756
rect 23852 18698 23863 18750
rect 23915 18698 23921 18750
rect 23852 16044 23908 18698
rect 23951 16265 24064 18820
rect 23945 16152 23951 16265
rect 24064 16152 24070 16265
rect 23852 15982 23908 15988
rect 23438 12790 23444 12846
rect 23500 12790 23506 12846
rect 23352 12784 23408 12790
rect 23260 11015 23316 12547
rect 23444 11808 23500 12790
rect 23444 11595 23500 11752
rect 23536 11680 23592 15548
rect 23951 15669 24064 15675
rect 24064 15625 24068 15631
rect 24064 15567 24068 15573
rect 23852 15486 23908 15492
rect 23852 15434 23863 15486
rect 23915 15434 23921 15486
rect 23852 12780 23908 15434
rect 23951 13001 24064 15556
rect 23945 12888 23951 13001
rect 24064 12888 24070 13001
rect 23852 12718 23908 12724
rect 23534 11674 23592 11680
rect 23586 11622 23592 11674
rect 23534 11616 23592 11622
rect 23536 11597 23592 11616
rect 23260 10953 23316 10959
rect 26888 10053 26946 12072
rect 26888 9989 26946 9995
rect 27164 9924 27222 12092
rect 27164 9860 27222 9866
rect 27439 9775 27497 12109
rect 27439 9711 27497 9717
rect 27714 9603 27772 12109
rect 27714 9539 27772 9545
rect 28271 9435 28329 12076
rect 28271 9371 28329 9377
rect 28391 9335 28449 12096
rect 28391 9271 28449 9277
rect 28511 9208 28569 12086
rect 28511 9144 28569 9150
rect 28631 9095 28689 12066
rect 28631 9031 28689 9037
<< metal4 >>
rect 56 35872 28639 40167
rect 56 23504 4351 35872
rect 18117 35472 22412 35872
rect 24344 35472 28639 35872
rect 13672 4311 17967 11984
rect 28789 4311 33084 11984
rect 8796 16 33084 4311
use SSTL  SSTL_0 ~/proj/caravan-project/mag/SSTL
timestamp 1644865263
transform 1 0 2350 0 -1 4308
box -2332 -19196 6668 4292
use SSTL  SSTL_1
timestamp 1644865263
transform -1 0 20118 0 -1 16276
box -2332 -19196 6668 4292
use SSTL  SSTL_2
timestamp 1644865263
transform 1 0 26638 0 -1 16276
box -2332 -19196 6668 4292
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform -1 0 23608 0 1 12576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1644111581
transform -1 0 23608 0 -1 15840
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1644111581
transform -1 0 23608 0 -1 19104
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1644111581
transform -1 0 23608 0 1 15840
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1644111581
transform -1 0 23608 0 -1 22368
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1644111581
transform -1 0 23608 0 1 19104
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1644111581
transform -1 0 23608 0 -1 25632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_7
timestamp 1644111581
transform -1 0 23608 0 1 22368
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_8
timestamp 1644111581
transform -1 0 23608 0 -1 28896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_9
timestamp 1644111581
transform -1 0 23608 0 1 25632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_10
timestamp 1644111581
transform -1 0 23608 0 -1 32160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_11
timestamp 1644111581
transform -1 0 23608 0 1 28896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_12
timestamp 1644111581
transform -1 0 23608 0 -1 35424
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_13
timestamp 1644111581
transform -1 0 23608 0 1 32160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 9716 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_1
timestamp 1644111581
transform 1 0 10084 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 12384 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 10452 0 1 11488
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 12752 0 1 11488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1644111581
transform 1 0 23608 0 1 12576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1644111581
transform 1 0 23608 0 -1 15840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1644111581
transform 1 0 23608 0 -1 19104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1644111581
transform 1 0 23608 0 1 15840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1644111581
transform 1 0 23608 0 -1 22368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1644111581
transform 1 0 23608 0 1 19104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1644111581
transform 1 0 23608 0 -1 25632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1644111581
transform 1 0 23608 0 1 22368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1644111581
transform 1 0 23608 0 -1 28896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1644111581
transform 1 0 23608 0 1 25632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1644111581
transform 1 0 23608 0 -1 32160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1644111581
transform 1 0 23608 0 1 28896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1644111581
transform 1 0 23608 0 -1 35424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1644111581
transform 1 0 23608 0 1 32160
box -38 -48 130 592
<< labels >>
flabel metal2 -276 16 -217 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[0]
port 8 n
flabel metal2 -156 16 -97 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[1]
port 9 n
flabel metal2 -36 16 23 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[2]
port 10 n
flabel metal2 84 16 143 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[3]
port 11 n
flabel metal2 204 16 263 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[4]
port 12 n
flabel metal2 324 16 383 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[5]
port 13 n
flabel metal2 444 16 503 112 1 FreeSerif 112 45 0 0 rx_leg_ctrl[6]
port 14 n
flabel metal2 2600 16 2658 112 1 FreeSerif 112 45 0 0 rx_pu_cal[0]
port 15 n
flabel metal2 2876 16 2934 112 1 FreeSerif 112 45 0 0 rx_pu_cal[1]
port 16 n
flabel metal2 3151 16 3209 112 1 FreeSerif 112 45 0 0 rx_pu_cal[2]
port 17 n
flabel metal2 3426 16 3484 112 1 FreeSerif 112 45 0 0 rx_pu_cal[3]
port 18 n
flabel metal2 3983 16 4041 112 1 FreeSerif 112 45 0 0 rx_pd_cal[0]
port 19 n
flabel metal2 4103 16 4161 112 1 FreeSerif 112 45 0 0 rx_pd_cal[1]
port 20 n
flabel metal2 4223 16 4281 112 1 FreeSerif 112 45 0 0 rx_pd_cal[2]
port 21 n
flabel metal2 4343 16 4401 112 1 FreeSerif 112 45 0 0 rx_pd_cal[3]
port 22 n
flabel metal2 6046 22576 6142 23504 1 FreeSerif 1600 0 0 0 rx_DQ
port 38 n
flabel metal2 30334 34175 30423 35472 1 FreeSerif 1600 0 0 0 tx_DQ
port 39 n
flabel metal2 16333 34122 16422 35472 1 FreeSerif 1600 0 0 0 n_tx_DQ
port 40 n
flabel metal2 s 11105 16 11165 108 1 FreeSerif 112 0 0 0 d_sel_0
port 1 n
flabel metal2 s 11663 16 11723 108 1 FreeSerif 112 0 0 0 d_sel_1
port 2 n
flabel metal2 s 10626 16 10700 108 1 FreeSerif 112 0 0 0 data_0
port 5 n
flabel metal2 s 10741 16 10773 108 1 FreeSerif 112 0 0 0 data_2
port 6 n
flabel metal2 s 10811 16 10860 108 1 FreeSerif 112 0 0 0 data_3
port 7 n
flabel metal2 s 18067 16 18125 108 1 FreeSerif 112 45 0 0 tx_pd_cal[3]
port 23 n
flabel metal2 s 18187 16 18245 108 1 FreeSerif 112 45 0 0 tx_pd_cal[2]
port 24 n
flabel metal2 s 18307 16 18365 108 1 FreeSerif 112 45 0 0 tx_pd_cal[1]
port 25 n
flabel metal2 s 18427 16 18485 108 1 FreeSerif 112 45 0 0 tx_pd_cal[0]
port 26 n
flabel metal2 s 18984 16 19042 108 1 FreeSerif 112 45 0 0 tx_pu_cal[3]
port 27 n
flabel metal2 s 19259 16 19317 108 1 FreeSerif 112 45 0 0 tx_pu_cal[2]
port 28 n
flabel metal2 s 19534 16 19592 108 1 FreeSerif 112 45 0 0 tx_pu_cal[1]
port 29 n
flabel metal2 s 19810 16 19868 108 1 FreeSerif 112 45 0 0 tx_pu_cal[0]
port 30 n
flabel metal2 s 22524 16 22580 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[0]
port 31 n
flabel metal2 s 22616 16 22672 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[1]
port 32 n
flabel metal2 s 22708 16 22764 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[2]
port 33 n
flabel metal2 s 22800 16 22856 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[3]
port 34 n
flabel metal2 s 22892 16 22948 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[4]
port 35 n
flabel metal2 s 22984 16 23040 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[5]
port 36 n
flabel metal2 s 23076 16 23132 108 1 FreeSerif 112 45 0 0 tx_leg_ctrl[6]
port 37 n
flabel metal4 56 35872 28639 40167 1 FreeSerif 4800 0 0 0 IO_VDD
port 41 n
flabel metal4 28789 16 33084 11984 1 FreeSerif 4800 0 0 0 IO_GND
port 42 n
flabel metal2 s 11890 16 11946 108 1 FreeSerif 112 0 0 0 dig_VDD
port 3 n
flabel metal2 s 12057 16 12113 108 1 FreeSerif 112 0 0 0 dig_GND
port 4 n
<< end >>
