magic
tech sky130A
magscale 1 2
timestamp 1646843053
<< error_p >>
rect -125 -65 -63 65
rect -33 -65 33 65
rect 63 -65 125 65
rect 155 -65 221 65
rect 251 -65 313 65
rect 343 -65 409 65
rect 439 -65 501 65
rect 531 -65 597 65
rect 627 -65 689 65
rect 719 -65 785 65
rect 815 -65 877 65
rect 907 -65 973 65
rect 1003 -65 1065 65
rect 1095 -65 1161 65
rect 1191 -65 1253 65
rect 1283 -65 1349 65
rect 1379 -65 1441 65
rect 1471 -65 1537 65
rect 1567 -65 1629 65
rect 1659 -65 1725 65
rect 1755 -65 1817 65
rect 1847 -65 1913 65
rect 1943 -65 2005 65
rect 2035 -65 2101 65
rect 2131 -65 2193 65
rect 2223 -65 2289 65
rect 2319 -65 2381 65
rect 2411 -65 2477 65
rect 2507 -65 2569 65
rect 2599 -65 2665 65
rect 2695 -65 2757 65
rect 2787 -65 2853 65
rect 2883 -65 2945 65
<< nmos >>
rect -63 -65 -33 65
rect 33 -65 63 65
rect 125 -65 155 65
rect 221 -65 251 65
rect 313 -65 343 65
rect 409 -65 439 65
rect 501 -65 531 65
rect 597 -65 627 65
rect 689 -65 719 65
rect 785 -65 815 65
rect 877 -65 907 65
rect 973 -65 1003 65
rect 1065 -65 1095 65
rect 1161 -65 1191 65
rect 1253 -65 1283 65
rect 1349 -65 1379 65
rect 1441 -65 1471 65
rect 1537 -65 1567 65
rect 1629 -65 1659 65
rect 1725 -65 1755 65
rect 1817 -65 1847 65
rect 1913 -65 1943 65
rect 2005 -65 2035 65
rect 2101 -65 2131 65
rect 2193 -65 2223 65
rect 2289 -65 2319 65
rect 2381 -65 2411 65
rect 2477 -65 2507 65
rect 2569 -65 2599 65
rect 2665 -65 2695 65
rect 2757 -65 2787 65
rect 2853 -65 2883 65
<< ndiff >>
rect -125 -17 -63 65
rect -125 -57 -113 -17
rect -79 -57 -63 -17
rect -125 -65 -63 -57
rect -33 57 33 65
rect -33 17 -17 57
rect 17 17 33 57
rect -33 -65 33 17
rect 63 -17 125 65
rect 63 -57 75 -17
rect 109 -57 125 -17
rect 63 -65 125 -57
rect 155 57 221 65
rect 155 17 171 57
rect 205 17 221 57
rect 155 -65 221 17
rect 251 -17 313 65
rect 251 -57 263 -17
rect 297 -57 313 -17
rect 251 -65 313 -57
rect 343 57 409 65
rect 343 17 359 57
rect 393 17 409 57
rect 343 -65 409 17
rect 439 -17 501 65
rect 439 -57 451 -17
rect 485 -57 501 -17
rect 439 -65 501 -57
rect 531 57 597 65
rect 531 17 547 57
rect 581 17 597 57
rect 531 -65 597 17
rect 627 -17 689 65
rect 627 -57 639 -17
rect 673 -57 689 -17
rect 627 -65 689 -57
rect 719 57 785 65
rect 719 17 735 57
rect 769 17 785 57
rect 719 -65 785 17
rect 815 -17 877 65
rect 815 -57 827 -17
rect 861 -57 877 -17
rect 815 -65 877 -57
rect 907 57 973 65
rect 907 17 923 57
rect 957 17 973 57
rect 907 -65 973 17
rect 1003 -17 1065 65
rect 1003 -57 1015 -17
rect 1049 -57 1065 -17
rect 1003 -65 1065 -57
rect 1095 57 1161 65
rect 1095 17 1111 57
rect 1145 17 1161 57
rect 1095 -65 1161 17
rect 1191 -17 1253 65
rect 1191 -57 1203 -17
rect 1237 -57 1253 -17
rect 1191 -65 1253 -57
rect 1283 57 1349 65
rect 1283 17 1299 57
rect 1333 17 1349 57
rect 1283 -65 1349 17
rect 1379 -17 1441 65
rect 1379 -57 1391 -17
rect 1425 -57 1441 -17
rect 1379 -65 1441 -57
rect 1471 57 1537 65
rect 1471 17 1487 57
rect 1521 17 1537 57
rect 1471 -65 1537 17
rect 1567 -17 1629 65
rect 1567 -57 1579 -17
rect 1613 -57 1629 -17
rect 1567 -65 1629 -57
rect 1659 57 1725 65
rect 1659 17 1675 57
rect 1709 17 1725 57
rect 1659 -65 1725 17
rect 1755 -17 1817 65
rect 1755 -57 1767 -17
rect 1801 -57 1817 -17
rect 1755 -65 1817 -57
rect 1847 57 1913 65
rect 1847 17 1863 57
rect 1897 17 1913 57
rect 1847 -65 1913 17
rect 1943 -17 2005 65
rect 1943 -57 1955 -17
rect 1989 -57 2005 -17
rect 1943 -65 2005 -57
rect 2035 57 2101 65
rect 2035 17 2051 57
rect 2085 17 2101 57
rect 2035 -65 2101 17
rect 2131 -17 2193 65
rect 2131 -57 2143 -17
rect 2177 -57 2193 -17
rect 2131 -65 2193 -57
rect 2223 57 2289 65
rect 2223 17 2239 57
rect 2273 17 2289 57
rect 2223 -65 2289 17
rect 2319 -17 2381 65
rect 2319 -57 2331 -17
rect 2365 -57 2381 -17
rect 2319 -65 2381 -57
rect 2411 57 2477 65
rect 2411 17 2427 57
rect 2461 17 2477 57
rect 2411 -65 2477 17
rect 2507 -17 2569 65
rect 2507 -57 2519 -17
rect 2553 -57 2569 -17
rect 2507 -65 2569 -57
rect 2599 57 2665 65
rect 2599 17 2615 57
rect 2649 17 2665 57
rect 2599 -65 2665 17
rect 2695 -17 2757 65
rect 2695 -57 2707 -17
rect 2741 -57 2757 -17
rect 2695 -65 2757 -57
rect 2787 57 2853 65
rect 2787 17 2803 57
rect 2837 17 2853 57
rect 2787 -65 2853 17
rect 2883 -17 2945 65
rect 2883 -57 2895 -17
rect 2929 -57 2945 -17
rect 2883 -65 2945 -57
<< ndiffc >>
rect -113 -57 -79 -17
rect -17 17 17 57
rect 75 -57 109 -17
rect 171 17 205 57
rect 263 -57 297 -17
rect 359 17 393 57
rect 451 -57 485 -17
rect 547 17 581 57
rect 639 -57 673 -17
rect 735 17 769 57
rect 827 -57 861 -17
rect 923 17 957 57
rect 1015 -57 1049 -17
rect 1111 17 1145 57
rect 1203 -57 1237 -17
rect 1299 17 1333 57
rect 1391 -57 1425 -17
rect 1487 17 1521 57
rect 1579 -57 1613 -17
rect 1675 17 1709 57
rect 1767 -57 1801 -17
rect 1863 17 1897 57
rect 1955 -57 1989 -17
rect 2051 17 2085 57
rect 2143 -57 2177 -17
rect 2239 17 2273 57
rect 2331 -57 2365 -17
rect 2427 17 2461 57
rect 2519 -57 2553 -17
rect 2615 17 2649 57
rect 2707 -57 2741 -17
rect 2803 17 2837 57
rect 2895 -57 2929 -17
<< poly >>
rect -63 65 -33 91
rect 33 65 63 91
rect 125 65 155 91
rect 221 65 251 91
rect 313 65 343 91
rect 409 65 439 91
rect 501 65 531 91
rect 597 65 627 91
rect 689 65 719 91
rect 785 65 815 91
rect 877 65 907 91
rect 973 65 1003 91
rect 1065 65 1095 91
rect 1161 65 1191 91
rect 1253 65 1283 91
rect 1349 65 1379 91
rect 1441 65 1471 91
rect 1537 65 1567 91
rect 1629 65 1659 91
rect 1725 65 1755 91
rect 1817 65 1847 91
rect 1913 65 1943 91
rect 2005 65 2035 91
rect 2101 65 2131 91
rect 2193 65 2223 91
rect 2289 65 2319 91
rect 2381 65 2411 91
rect 2477 65 2507 91
rect 2569 65 2599 91
rect 2665 65 2695 91
rect 2757 65 2787 91
rect 2853 65 2883 91
rect -63 -87 -33 -65
rect 33 -87 63 -65
rect 125 -87 155 -65
rect 221 -87 251 -65
rect 313 -87 343 -65
rect 409 -87 439 -65
rect 501 -87 531 -65
rect 597 -87 627 -65
rect 689 -87 719 -65
rect 785 -87 815 -65
rect 877 -87 907 -65
rect 973 -87 1003 -65
rect 1065 -87 1095 -65
rect 1161 -87 1191 -65
rect 1253 -87 1283 -65
rect 1349 -87 1379 -65
rect 1441 -87 1471 -65
rect 1537 -87 1567 -65
rect 1629 -87 1659 -65
rect 1725 -87 1755 -65
rect 1817 -87 1847 -65
rect 1913 -87 1943 -65
rect 2005 -87 2035 -65
rect 2101 -87 2131 -65
rect 2193 -87 2223 -65
rect 2289 -87 2319 -65
rect 2381 -87 2411 -65
rect 2477 -87 2507 -65
rect 2569 -87 2599 -65
rect 2665 -87 2695 -65
rect 2757 -87 2787 -65
rect 2853 -87 2883 -65
rect -125 -103 2901 -87
rect -125 -137 -65 -103
rect -31 -137 31 -103
rect 65 -137 123 -103
rect 157 -137 219 -103
rect 253 -137 311 -103
rect 345 -137 407 -103
rect 441 -137 499 -103
rect 533 -137 595 -103
rect 629 -137 687 -103
rect 721 -137 783 -103
rect 817 -137 875 -103
rect 909 -137 971 -103
rect 1005 -137 1063 -103
rect 1097 -137 1159 -103
rect 1193 -137 1251 -103
rect 1285 -137 1347 -103
rect 1381 -137 1439 -103
rect 1473 -137 1535 -103
rect 1569 -137 1627 -103
rect 1661 -137 1723 -103
rect 1757 -137 1815 -103
rect 1849 -137 1911 -103
rect 1945 -137 2003 -103
rect 2037 -137 2099 -103
rect 2133 -137 2191 -103
rect 2225 -137 2287 -103
rect 2321 -137 2379 -103
rect 2413 -137 2475 -103
rect 2509 -137 2567 -103
rect 2601 -137 2663 -103
rect 2697 -137 2755 -103
rect 2789 -137 2851 -103
rect 2885 -137 2901 -103
rect -125 -153 2901 -137
<< polycont >>
rect -65 -137 -31 -103
rect 31 -137 65 -103
rect 123 -137 157 -103
rect 219 -137 253 -103
rect 311 -137 345 -103
rect 407 -137 441 -103
rect 499 -137 533 -103
rect 595 -137 629 -103
rect 687 -137 721 -103
rect 783 -137 817 -103
rect 875 -137 909 -103
rect 971 -137 1005 -103
rect 1063 -137 1097 -103
rect 1159 -137 1193 -103
rect 1251 -137 1285 -103
rect 1347 -137 1381 -103
rect 1439 -137 1473 -103
rect 1535 -137 1569 -103
rect 1627 -137 1661 -103
rect 1723 -137 1757 -103
rect 1815 -137 1849 -103
rect 1911 -137 1945 -103
rect 2003 -137 2037 -103
rect 2099 -137 2133 -103
rect 2191 -137 2225 -103
rect 2287 -137 2321 -103
rect 2379 -137 2413 -103
rect 2475 -137 2509 -103
rect 2567 -137 2601 -103
rect 2663 -137 2697 -103
rect 2755 -137 2789 -103
rect 2851 -137 2885 -103
<< locali >>
rect -125 17 -17 57
rect 17 17 171 57
rect 205 17 359 57
rect 393 17 547 57
rect 581 17 735 57
rect 769 17 923 57
rect 957 17 1111 57
rect 1145 17 1299 57
rect 1333 17 1487 57
rect 1521 17 1675 57
rect 1709 17 1863 57
rect 1897 17 2051 57
rect 2085 17 2239 57
rect 2273 17 2427 57
rect 2461 17 2615 57
rect 2649 17 2803 57
rect 2837 17 2945 57
rect -129 -57 -113 -17
rect -79 -57 75 -17
rect 109 -57 263 -17
rect 297 -57 451 -17
rect 485 -57 639 -17
rect 673 -57 827 -17
rect 861 -57 1015 -17
rect 1049 -57 1203 -17
rect 1237 -57 1391 -17
rect 1425 -57 1579 -17
rect 1613 -57 1767 -17
rect 1801 -57 1955 -17
rect 1989 -57 2143 -17
rect 2177 -57 2331 -17
rect 2365 -57 2519 -17
rect 2553 -57 2707 -17
rect 2741 -57 2895 -17
rect 2929 -57 2945 -17
rect -125 -137 -65 -103
rect -31 -137 31 -103
rect 65 -137 123 -103
rect 157 -137 219 -103
rect 253 -137 311 -103
rect 345 -137 407 -103
rect 441 -137 499 -103
rect 533 -137 595 -103
rect 629 -137 687 -103
rect 721 -137 783 -103
rect 817 -137 875 -103
rect 909 -137 971 -103
rect 1005 -137 1063 -103
rect 1097 -137 1159 -103
rect 1193 -137 1251 -103
rect 1285 -137 1347 -103
rect 1381 -137 1439 -103
rect 1473 -137 1535 -103
rect 1569 -137 1627 -103
rect 1661 -137 1723 -103
rect 1757 -137 1815 -103
rect 1849 -137 1911 -103
rect 1945 -137 2003 -103
rect 2037 -137 2099 -103
rect 2133 -137 2191 -103
rect 2225 -137 2287 -103
rect 2321 -137 2379 -103
rect 2413 -137 2475 -103
rect 2509 -137 2567 -103
rect 2601 -137 2663 -103
rect 2697 -137 2755 -103
rect 2789 -137 2851 -103
rect 2885 -137 2901 -103
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.650 l 0.150 m 1 nf 2 diffcov 25 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
