* NGSPICE file created from SSTL.ext - technology: sky130A

.subckt n-leg_ctrl_fet_2 a_n125_n65# a_n81_n153# a_n33_n65# VSUBS
X0 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=4.03e+11p ps=3.84e+06u w=650000u l=150000u
X1 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n125_n65# a_n81_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_n81_n153# a_n125_n65# 0.13fF
C1 a_n81_n153# a_n33_n65# 0.24fF
C2 a_n125_n65# a_n33_n65# 0.45fF
C3 a_n33_n65# VSUBS 0.02fF
C4 a_n125_n65# VSUBS 0.02fF
C5 a_n81_n153# VSUBS 0.33fF
.ends

.subckt n-leg_ctrl_fet_0 a_n125_n153# a_n125_n65# a_n33_n65# VSUBS
X0 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=3.4255e+12p pd=3.264e+07u as=3.432e+12p ps=3.136e+07u w=650000u l=150000u
X1 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_n33_n65# a_n125_n153# 1.42fF
C1 a_n33_n65# a_n125_n65# 3.92fF
C2 a_n125_n65# a_n125_n153# 2.76fF
C3 a_n33_n65# VSUBS 0.02fF
C4 a_n125_n65# VSUBS 0.02fF
C5 a_n125_n153# VSUBS 3.21fF
.ends

.subckt n-leg_ctrl_fet_3 a_15_n19# a_n73_n19# a_n33_n107# VSUBS
X0 a_15_n19# a_n33_n107# a_n73_n19# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
C0 a_15_n19# a_n73_n19# 0.07fF
C1 a_15_n19# VSUBS 0.02fF
C2 a_n73_n19# VSUBS 0.02fF
C3 a_n33_n107# VSUBS 0.13fF
.ends

.subckt n-leg_ctrl_fet_1 a_n125_n153# a_n125_n65# a_n33_n65# VSUBS
X0 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=7.84e+06u as=1.0075e+12p ps=9.6e+06u w=650000u l=150000u
X1 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_n125_n65# a_n33_n65# 1.05fF
C1 a_n125_n65# a_n125_n153# 0.37fF
C2 a_n125_n153# a_n33_n65# 0.73fF
C3 a_n33_n65# VSUBS 0.02fF
C4 a_n125_n65# VSUBS 0.02fF
C5 a_n125_n153# VSUBS 0.88fF
.ends

.subckt n-leg_polyres a_n33_170# a_n33_n243# VSUBS
R0 a_n33_n243# a_n33_170# sky130_fd_pr__res_generic_po w=330000u l=1.7e+06u
C0 a_n33_170# a_n33_n243# 0.01fF
C1 a_n33_n243# VSUBS 0.07fF
C2 a_n33_170# VSUBS 0.07fF
.ends

.subckt n-leg pd_ctrl cal_ctrl[0] cal_ctrl[1] cal_ctrl[2] cal_ctrl[3] li_1854_527#
+ vpulldown DQ GND
Xn-leg_ctrl_fet_2_0 DQ cal_ctrl[2] vpulldown GND n-leg_ctrl_fet_2
Xn-leg_ctrl_fet_0_0 cal_ctrl[0] DQ vpulldown GND n-leg_ctrl_fet_0
Xn-leg_ctrl_fet_3_0 DQ vpulldown cal_ctrl[3] GND n-leg_ctrl_fet_3
Xn-leg_ctrl_fet_1_0 cal_ctrl[1] vpulldown DQ GND n-leg_ctrl_fet_1
Xn-leg_polyres_0 vpulldown DQ GND n-leg_polyres
X0 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=1.20215e+13p pd=2.595e+06u as=9.6163e+12p ps=9.0425e+07u w=650000u l=150000u
X1 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X42 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 cal_ctrl[2] DQ 0.26fF
C1 li_1854_527# cal_ctrl[0] 0.56fF
C2 cal_ctrl[0] cal_ctrl[3] 0.73fF
C3 li_1854_527# cal_ctrl[3] 5.59fF
C4 vpulldown cal_ctrl[1] 0.76fF
C5 pd_ctrl vpulldown 7.80fF
C6 cal_ctrl[0] cal_ctrl[2] 0.98fF
C7 li_1854_527# cal_ctrl[2] 1.94fF
C8 cal_ctrl[2] cal_ctrl[3] 7.56fF
C9 DQ cal_ctrl[1] 1.18fF
C10 pd_ctrl DQ 0.03fF
C11 vpulldown DQ 0.55fF
C12 cal_ctrl[0] cal_ctrl[1] 5.93fF
C13 li_1854_527# cal_ctrl[1] 0.87fF
C14 cal_ctrl[3] cal_ctrl[1] 1.18fF
C15 li_1854_527# pd_ctrl 0.55fF
C16 cal_ctrl[0] vpulldown 0.08fF
C17 li_1854_527# vpulldown 2.00fF
C18 vpulldown cal_ctrl[3] 0.17fF
C19 cal_ctrl[2] cal_ctrl[1] 2.56fF
C20 cal_ctrl[0] DQ 0.18fF
C21 cal_ctrl[2] vpulldown 0.86fF
C22 li_1854_527# DQ 0.80fF
C23 DQ cal_ctrl[3] 0.15fF
C24 pd_ctrl GND 8.51fF
C25 li_1854_527# GND 4.28fF
C26 DQ GND 1.52fF
C27 vpulldown GND 12.60fF
C28 cal_ctrl[1] GND 4.42fF
C29 cal_ctrl[3] GND 2.77fF
C30 cal_ctrl[0] GND 13.30fF
C31 cal_ctrl[2] GND 2.75fF
.ends

.subckt p-leg_fet_16 a_n1053_n161# a_n1053_n64# a_995_n64# a_n285_n64# a_n541_n64#
+ a_483_n64# a_739_n64# a_n29_n64# a_n925_n64# a_227_n64# w_n1089_n100# a_n797_n64#
+ VSUBS
X0 a_n925_n64# a_n1053_n161# a_n541_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n797_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X2 a_n925_n64# a_n1053_n161# a_227_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X3 a_739_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X4 a_n925_n64# a_n1053_n161# a_n29_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_n285_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X6 a_n925_n64# a_n1053_n161# a_n797_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X7 a_227_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X8 a_n925_n64# a_n1053_n161# a_483_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X9 a_995_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X10 a_n925_n64# a_n1053_n161# a_n1053_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X11 a_n925_n64# a_n1053_n161# a_739_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X12 a_n541_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X13 a_n925_n64# a_n1053_n161# a_n285_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X14 a_n29_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X15 a_483_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
C0 a_n541_n64# a_n797_n64# 0.02fF
C1 a_227_n64# a_n925_n64# 0.06fF
C2 a_995_n64# w_n1089_n100# 0.07fF
C3 a_n925_n64# a_n1053_n64# 0.07fF
C4 a_227_n64# a_n29_n64# 0.02fF
C5 a_227_n64# a_483_n64# 0.02fF
C6 a_n797_n64# w_n1089_n100# 0.07fF
C7 a_739_n64# w_n1089_n100# 0.07fF
C8 a_n925_n64# a_n1053_n161# 2.38fF
C9 a_739_n64# a_995_n64# 0.02fF
C10 a_n29_n64# a_n925_n64# 0.06fF
C11 a_n925_n64# a_483_n64# 0.06fF
C12 a_n925_n64# a_n285_n64# 0.06fF
C13 a_n925_n64# a_n541_n64# 0.06fF
C14 a_227_n64# w_n1089_n100# 0.07fF
C15 a_n29_n64# a_n285_n64# 0.02fF
C16 a_n1053_n64# w_n1089_n100# 0.07fF
C17 a_n541_n64# a_n285_n64# 0.02fF
C18 a_n925_n64# w_n1089_n100# 1.05fF
C19 a_n925_n64# a_995_n64# 0.07fF
C20 a_n1053_n161# w_n1089_n100# 0.95fF
C21 a_n29_n64# w_n1089_n100# 0.07fF
C22 a_483_n64# w_n1089_n100# 0.07fF
C23 a_n797_n64# a_n1053_n64# 0.02fF
C24 a_n285_n64# w_n1089_n100# 0.07fF
C25 a_n541_n64# w_n1089_n100# 0.07fF
C26 a_n925_n64# a_n797_n64# 0.06fF
C27 a_n925_n64# a_739_n64# 0.06fF
C28 a_483_n64# a_739_n64# 0.02fF
C29 a_995_n64# VSUBS -0.04fF
C30 a_739_n64# VSUBS -0.04fF
C31 a_483_n64# VSUBS -0.04fF
C32 a_227_n64# VSUBS -0.04fF
C33 a_n29_n64# VSUBS -0.04fF
C34 a_n285_n64# VSUBS -0.04fF
C35 a_n541_n64# VSUBS -0.04fF
C36 a_n797_n64# VSUBS -0.04fF
C37 a_n925_n64# VSUBS -0.84fF
C38 a_n1053_n64# VSUBS -0.04fF
C39 a_n1053_n161# VSUBS 1.21fF
C40 w_n1089_n100# VSUBS 1.95fF
.ends

.subckt p-leg_polyres a_n33_n253# a_n33_180# VSUBS
R0 a_n33_n253# a_n33_180# sky130_fd_pr__res_generic_po w=330000u l=1.8e+06u
C0 a_n33_n253# VSUBS 0.09fF
C1 a_n33_180# VSUBS 0.09fF
.ends

.subckt p-leg_6 a_n1053_n64# a_n285_n64# a_n541_n64# a_n995_n161# a_n925_n64# w_n1089_n100#
+ a_n797_n64# VSUBS
X0 a_n925_n64# a_n995_n161# a_n541_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n797_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X2 a_n285_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X3 a_n925_n64# a_n995_n161# a_n797_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4 a_n925_n64# a_n995_n161# a_n1053_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_n541_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
C0 a_n925_n64# a_n797_n64# 0.06fF
C1 a_n541_n64# a_n797_n64# 0.02fF
C2 w_n1089_n100# a_n797_n64# 0.06fF
C3 a_n925_n64# a_n541_n64# 0.06fF
C4 a_n925_n64# w_n1089_n100# 0.42fF
C5 a_n925_n64# a_n995_n161# 0.84fF
C6 a_n541_n64# w_n1089_n100# 0.06fF
C7 a_n995_n161# w_n1089_n100# 0.34fF
C8 a_n925_n64# a_n285_n64# 0.06fF
C9 a_n541_n64# a_n285_n64# 0.02fF
C10 a_n1053_n64# a_n797_n64# 0.02fF
C11 w_n1089_n100# a_n285_n64# 0.06fF
C12 a_n925_n64# a_n1053_n64# 0.07fF
C13 a_n1053_n64# w_n1089_n100# 0.06fF
C14 a_n285_n64# VSUBS -0.05fF
C15 a_n541_n64# VSUBS -0.05fF
C16 a_n797_n64# VSUBS -0.05fF
C17 a_n925_n64# VSUBS -0.33fF
C18 a_n1053_n64# VSUBS -0.05fF
C19 a_n995_n161# VSUBS 0.44fF
C20 w_n1089_n100# VSUBS 0.80fF
.ends

.subckt p-leg n_cal_ctrl[0] n_cal_ctrl[1] n_cal_ctrl[2] n_cal_ctrl[3] w_3710_2162#
+ li_4_2169# w_1502_2162# w_4446_2162# w_2974_2162# w_2238_2162# w_5918_2162# extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ w_766_2162# extr_sky130_fd_sc_hd__fill_8_8/VGND extr_sky130_fd_sc_hd__fill_8_9/VGND VDD li_16_1957#
+ w_5182_2162# n_pu_ctrl p-leg_6_6/VSUBS DQ
Xp-leg_fet_16_4 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
Xp-leg_fet_16_5 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
Xp-leg_fet_16_6 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_6_6/VSUBS p-leg_fet_16
Xp-leg_fet_16_7 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_6_6/VSUBS p-leg_fet_16
Xp-leg_polyres_0 DQ li_16_1957# p-leg_6_6/VSUBS p-leg_polyres
Xp-leg_fet_16_8 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_6_6/VSUBS p-leg_fet_16
Xp-leg_6_0 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_6_1 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_6_2 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_6_3 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_6_4 DQ DQ DQ n_cal_ctrl[2] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_6_6 li_16_1957# li_16_1957# li_16_1957# n_cal_ctrl[3] DQ VDD li_16_1957# p-leg_6_6/VSUBS
+ p-leg_6
Xp-leg_6_5 DQ DQ DQ n_cal_ctrl[2] li_16_1957# VDD DQ p-leg_6_6/VSUBS p-leg_6
Xp-leg_fet_16_0 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
Xp-leg_fet_16_1 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
Xp-leg_fet_16_2 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
Xp-leg_fet_16_3 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_6_6/VSUBS
+ p-leg_fet_16
C0 extr_sky130_fd_sc_hd__fill_8_8/VGND VDD 0.08fF
C1 li_16_1957# VDD 5.24fF
C2 li_16_1957# n_cal_ctrl[2] 1.83fF
C3 n_pu_ctrl extr_sky130_fd_sc_hd__fill_8_8/VGND 1.13fF
C4 n_pu_ctrl li_16_1957# 0.03fF
C5 li_16_1957# n_cal_ctrl[3] 1.50fF
C6 li_16_1957# extr_sky130_fd_sc_hd__fill_8_9/VGND 1.97fF
C7 li_16_1957# n_cal_ctrl[0] 3.57fF
C8 li_16_1957# DQ 6.76fF
C9 extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C10 li_4_2169# n_cal_ctrl[0] 0.80fF
C11 li_4_2169# DQ 0.72fF
C12 n_cal_ctrl[2] VDD 6.76fF
C13 n_pu_ctrl VDD 2.31fF
C14 n_pu_ctrl n_cal_ctrl[2] 0.08fF
C15 li_16_1957# n_cal_ctrl[1] 1.06fF
C16 n_cal_ctrl[3] VDD 2.74fF
C17 extr_sky130_fd_sc_hd__fill_8_9/VGND VDD 0.34fF
C18 n_cal_ctrl[0] VDD 20.34fF
C19 n_cal_ctrl[3] n_cal_ctrl[2] 7.51fF
C20 n_cal_ctrl[2] extr_sky130_fd_sc_hd__fill_8_9/VGND 1.84fF
C21 DQ VDD 3.33fF
C22 n_cal_ctrl[2] n_cal_ctrl[0] 1.44fF
C23 n_pu_ctrl n_cal_ctrl[3] 0.14fF
C24 n_pu_ctrl extr_sky130_fd_sc_hd__fill_8_9/VGND 1.32fF
C25 n_cal_ctrl[2] DQ 2.44fF
C26 n_pu_ctrl DQ 0.59fF
C27 n_cal_ctrl[1] VDD 16.25fF
C28 n_cal_ctrl[2] n_cal_ctrl[1] 7.25fF
C29 n_cal_ctrl[3] extr_sky130_fd_sc_hd__fill_8_9/VGND 2.41fF
C30 n_pu_ctrl n_cal_ctrl[1] 0.12fF
C31 n_cal_ctrl[3] n_cal_ctrl[0] 0.52fF
C32 n_cal_ctrl[3] DQ 2.21fF
C33 DQ extr_sky130_fd_sc_hd__fill_8_9/VGND 2.25fF
C34 li_16_1957# extr_sky130_fd_sc_hd__fill_8_8/VGND 0.78fF
C35 DQ n_cal_ctrl[0] 0.53fF
C36 li_4_2169# li_16_1957# 2.07fF
C37 n_cal_ctrl[3] n_cal_ctrl[1] 2.02fF
C38 extr_sky130_fd_sc_hd__fill_8_9/VGND n_cal_ctrl[1] 0.80fF
C39 n_cal_ctrl[0] n_cal_ctrl[1] 3.06fF
C40 DQ n_cal_ctrl[1] 1.68fF
C41 n_cal_ctrl[1] p-leg_6_6/VSUBS -0.59fF
C42 li_4_2169# p-leg_6_6/VSUBS 6.04fF
C43 VDD p-leg_6_6/VSUBS 33.14fF
C44 n_cal_ctrl[3] p-leg_6_6/VSUBS 1.75fF
C45 extr_sky130_fd_sc_hd__fill_8_9/VPWR p-leg_6_6/VSUBS 0.16fF
C46 n_cal_ctrl[2] p-leg_6_6/VSUBS -0.44fF
C47 DQ p-leg_6_6/VSUBS -3.95fF
C48 li_16_1957# p-leg_6_6/VSUBS -6.69fF
C49 extr_sky130_fd_sc_hd__fill_8_8/VGND p-leg_6_6/VSUBS 6.12fF
C50 n_cal_ctrl[0] p-leg_6_6/VSUBS 0.18fF
C51 extr_sky130_fd_sc_hd__fill_8_9/VGND p-leg_6_6/VSUBS 5.24fF
C52 n_pu_ctrl p-leg_6_6/VSUBS 6.68fF
.ends

.subckt extr_sky130_fd_sc_hd__clkbuf_8 A VGND VPWR X a_110_47# VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=6.951e+11p ps=8.35e+06u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPWR VPB 1.16fF
C1 VPWR A 0.08fF
C2 X a_110_47# 1.39fF
C3 X VPB 0.51fF
C4 X VPWR 1.77fF
C5 VGND a_110_47# 0.43fF
C6 VGND A 0.08fF
C7 VGND VPWR 0.05fF
C8 a_110_47# VPB 0.65fF
C9 a_110_47# A 0.39fF
C10 VPWR a_110_47# 0.68fF
C11 VGND X 1.10fF
C12 VPB A 0.12fF
C13 VGND VNB 0.81fF
C14 X VNB -0.20fF
C15 VPWR VNB -0.38fF
C16 A VNB 0.34fF
C17 VPB VNB 1.05fF
C18 a_110_47# VNB 0.94fF
.ends

.subckt extr_sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VGND Y 0.67fF
C1 VPWR A 0.16fF
C2 VPB A 0.25fF
C3 VPWR VPB 0.76fF
C4 VGND A 0.16fF
C5 VPWR VGND 0.02fF
C6 Y A 1.17fF
C7 VPWR Y 1.39fF
C8 VPB Y 0.47fF
C9 VGND VNB 0.55fF
C10 Y VNB -0.02fF
C11 VPWR VNB -0.25fF
C12 A VNB 0.70fF
C13 VPB VNB 0.69fF
.ends

.subckt extr_sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 A VGND 0.87fF
C1 VPB Y 1.61fF
C2 VPWR Y 4.93fF
C3 VGND Y 1.83fF
C4 A Y 2.06fF
C5 VPWR VPB 2.42fF
C6 VPWR VGND 0.08fF
C7 VPB A 1.33fF
C8 VPWR A 0.81fF
C9 VGND VNB 1.80fF
C10 Y VNB -1.03fF
C11 VPWR VNB -0.94fF
C12 A VNB 2.35fF
C13 VPB VNB 2.20fF
.ends

.subckt extr_sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X a_110_47# VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPWR VPB 1.97fF
C1 a_110_47# VPB 1.36fF
C2 VPWR X 3.42fF
C3 VPWR VGND 0.07fF
C4 a_110_47# X 3.32fF
C5 A VPWR 0.08fF
C6 a_110_47# VGND 0.95fF
C7 A a_110_47# 0.54fF
C8 X VPB 1.02fF
C9 A VPB 0.21fF
C10 X VGND 2.23fF
C11 VPWR a_110_47# 1.15fF
C12 A VGND 0.12fF
C13 VGND VNB 1.41fF
C14 X VNB -0.49fF
C15 VPWR VNB -0.69fF
C16 A VNB 0.59fF
C17 VPB VNB 1.85fF
C18 a_110_47# VNB 1.82fF
.ends

.subckt extr_sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
C0 VPB Y 0.12fF
C1 Y VGND 0.20fF
C2 VPB A 0.07fF
C3 Y A 0.14fF
C4 VGND A 0.06fF
C5 VPB VPWR 0.33fF
C6 Y VPWR 0.26fF
C7 VGND VPWR 0.01fF
C8 A VPWR 0.06fF
C9 VGND VNB 0.37fF
C10 Y VNB 0.06fF
C11 VPWR VNB -0.02fF
C12 A VNB 0.15fF
C13 VPB VNB 0.34fF
.ends

.subckt SSTL DQ GND pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3] pd_ctrl[0]
+ pd_ctrl[1] pd_ctrl[2] pd_ctrl[3] pd_ctrl[4] pd_ctrl[5] pd_ctrl[6] pu_cal_ctrl[0]
+ pu_cal_ctrl[1] pu_cal_ctrl[2] pu_cal_ctrl[3] pu_ctrl[0] pu_ctrl[1] pu_ctrl[2] pu_ctrl[3]
+ pu_ctrl[4] pu_ctrl[5] pu_ctrl[6] VDD
Xn-leg_0 n-leg_0/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_0/vpulldown DQ GND n-leg
Xp-leg_3 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_3/w_3710_2162# GND p-leg_3/w_1502_2162# p-leg_3/w_4446_2162# p-leg_3/w_2974_2162#
+ p-leg_3/w_2238_2162# p-leg_3/w_5918_2162# p-leg_3/extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ p-leg_3/w_766_2162# GND GND VDD p-leg_3/li_16_1957# p-leg_3/w_5182_2162# p-leg_3/n_pu_ctrl
+ GND DQ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_1 extr_sky130_fd_sc_hd__clkinv_4_2/Y GND VDD n-leg_1/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xn-leg_1 n-leg_1/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_1/vpulldown DQ GND n-leg
Xp-leg_4 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_4/w_3710_2162# GND p-leg_4/w_1502_2162# p-leg_4/w_4446_2162# p-leg_4/w_2974_2162#
+ p-leg_4/w_2238_2162# p-leg_4/w_5918_2162# p-leg_4/extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ p-leg_4/w_766_2162# GND GND VDD p-leg_4/li_16_1957# p-leg_4/w_5182_2162# p-leg_4/n_pu_ctrl
+ GND DQ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_2 extr_sky130_fd_sc_hd__clkinv_4_4/Y GND VDD n-leg_2/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xn-leg_2 n-leg_2/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_2/vpulldown DQ GND n-leg
Xp-leg_5 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_5/w_3710_2162# GND p-leg_5/w_1502_2162# p-leg_5/w_4446_2162# p-leg_5/w_2974_2162#
+ p-leg_5/w_2238_2162# p-leg_5/w_5918_2162# VDD p-leg_5/w_766_2162# GND GND VDD p-leg_5/li_16_1957#
+ p-leg_5/w_5182_2162# p-leg_5/n_pu_ctrl GND DQ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_3 extr_sky130_fd_sc_hd__clkinv_4_6/Y GND VDD n-leg_3/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_10 extr_sky130_fd_sc_hd__clkinv_4_11/Y GND VDD extr_sky130_fd_sc_hd__clkbuf_8_5/A
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_3 n-leg_3/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_3/vpulldown DQ GND n-leg
Xp-leg_6 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_6/w_3710_2162# GND p-leg_6/w_1502_2162# p-leg_6/w_4446_2162# p-leg_6/w_2974_2162#
+ p-leg_6/w_2238_2162# p-leg_6/w_5918_2162# p-leg_6/extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ p-leg_6/w_766_2162# GND GND VDD p-leg_6/li_16_1957# p-leg_6/w_5182_2162# p-leg_6/n_pu_ctrl
+ GND DQ p-leg
Xextr_sky130_fd_sc_hd__clkinv_16_0 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_4 extr_sky130_fd_sc_hd__clkinv_4_8/Y GND VDD n-leg_4/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_11 pd_ctrl[5] GND VDD extr_sky130_fd_sc_hd__clkinv_4_11/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_4 n-leg_4/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_4/vpulldown DQ GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_16_1 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_5 extr_sky130_fd_sc_hd__clkbuf_8_5/A GND VDD n-leg_5/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_12 extr_sky130_fd_sc_hd__clkinv_4_13/Y GND VDD extr_sky130_fd_sc_hd__clkbuf_8_6/A
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_5 n-leg_5/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_5/vpulldown DQ GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_16_2 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_6 extr_sky130_fd_sc_hd__clkbuf_8_6/A GND VDD n-leg_6/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_13 pd_ctrl[6] GND VDD extr_sky130_fd_sc_hd__clkinv_4_13/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_6 n-leg_6/pd_ctrl pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD n-leg_6/vpulldown DQ GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_4_0 extr_sky130_fd_sc_hd__clkinv_4_1/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_0/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_3 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_1 pd_ctrl[0] GND VDD extr_sky130_fd_sc_hd__clkinv_4_1/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_4 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_2 extr_sky130_fd_sc_hd__clkinv_4_3/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_2/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_5 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_3 pd_ctrl[1] GND VDD extr_sky130_fd_sc_hd__clkinv_4_3/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_6 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_4 extr_sky130_fd_sc_hd__clkinv_4_5/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_4/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_7 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_5 pd_ctrl[2] GND VDD extr_sky130_fd_sc_hd__clkinv_4_5/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_8 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_20 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_6 extr_sky130_fd_sc_hd__clkinv_4_7/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_6/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_9 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_10 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_7 pd_ctrl[3] GND VDD extr_sky130_fd_sc_hd__clkinv_4_7/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_4_8 extr_sky130_fd_sc_hd__clkinv_4_9/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_8/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_11 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_12 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_9 pd_ctrl[4] GND VDD extr_sky130_fd_sc_hd__clkinv_4_9/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_13 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_14 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_15 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_16 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_0 pu_ctrl[0] GND VDD extr_sky130_fd_sc_hd__clkinv_16_2/A extr_sky130_fd_sc_hd__clkbuf_16_0/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_17 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_1 pu_ctrl[1] GND VDD extr_sky130_fd_sc_hd__clkinv_16_5/A extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_18 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_2 pu_ctrl[2] GND VDD extr_sky130_fd_sc_hd__clkinv_16_8/A extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_19 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_3 pu_ctrl[3] GND VDD extr_sky130_fd_sc_hd__clkinv_16_9/A extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_4 pu_ctrl[4] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_4/X extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_5 pu_ctrl[5] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_5/X extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_6 pu_ctrl[6] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_6/X extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47#
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__inv_1_0 pu_cal_ctrl[0] GND VDD p-leg_6/n_cal_ctrl[0] GND VDD extr_sky130_fd_sc_hd__inv_1
Xextr_sky130_fd_sc_hd__inv_1_1 pu_cal_ctrl[1] GND VDD p-leg_6/n_cal_ctrl[1] GND VDD extr_sky130_fd_sc_hd__inv_1
Xp-leg_0 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ GND GND GND GND GND GND GND p-leg_0/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND GND GND VDD
+ p-leg_0/li_16_1957# GND p-leg_0/n_pu_ctrl GND DQ p-leg
Xp-leg_1 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_1/w_3710_2162# GND p-leg_1/w_1502_2162# p-leg_1/w_4446_2162# p-leg_1/w_2974_2162#
+ p-leg_1/w_2238_2162# p-leg_1/w_5918_2162# p-leg_1/extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ p-leg_1/w_766_2162# GND GND VDD p-leg_1/li_16_1957# p-leg_1/w_5182_2162# p-leg_1/n_pu_ctrl
+ GND DQ p-leg
Xextr_sky130_fd_sc_hd__inv_1_2 pu_cal_ctrl[2] GND VDD p-leg_6/n_cal_ctrl[2] GND VDD extr_sky130_fd_sc_hd__inv_1
Xextr_sky130_fd_sc_hd__inv_1_3 pu_cal_ctrl[3] GND VDD p-leg_6/n_cal_ctrl[3] GND VDD extr_sky130_fd_sc_hd__inv_1
Xp-leg_2 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[3]
+ p-leg_2/w_3710_2162# GND p-leg_2/w_1502_2162# p-leg_2/w_4446_2162# p-leg_2/w_2974_2162#
+ p-leg_2/w_2238_2162# p-leg_2/w_5918_2162# VDD p-leg_2/w_766_2162# GND GND VDD p-leg_2/li_16_1957#
+ p-leg_2/w_5182_2162# p-leg_2/n_pu_ctrl GND DQ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_0 extr_sky130_fd_sc_hd__clkinv_4_0/Y GND VDD n-leg_0/pd_ctrl
+ extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# GND VDD extr_sky130_fd_sc_hd__clkbuf_8
C0 extr_sky130_fd_sc_hd__clkbuf_8_5/A extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.28fF
C1 extr_sky130_fd_sc_hd__clkbuf_8_6/A VDD 0.15fF
C2 extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_8/Y 0.05fF
C3 pd_cal_ctrl[3] p-leg_6/n_cal_ctrl[1] 1.62fF
C4 p-leg_4/li_16_1957# VDD 0.01fF
C5 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# VDD 0.05fF
C6 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C7 pd_cal_ctrl[3] p-leg_6/n_cal_ctrl[2] 0.45fF
C8 p-leg_2/li_16_1957# pd_cal_ctrl[0] 0.66fF
C9 extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_13/Y 0.01fF
C10 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# VDD 0.05fF
C11 pu_cal_ctrl[0] pu_cal_ctrl[1] 0.13fF
C12 extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.03fF
C13 p-leg_3/n_pu_ctrl p-leg_6/n_cal_ctrl[1] 0.35fF
C14 p-leg_2/li_16_1957# p-leg_2/n_pu_ctrl 0.30fF
C15 p-leg_0/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.39fF
C16 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[3] 1.67fF
C17 p-leg_6/n_cal_ctrl[0] p-leg_4/n_pu_ctrl 0.58fF
C18 VDD n-leg_5/pd_ctrl 0.06fF
C19 pd_cal_ctrl[0] p-leg_2/n_pu_ctrl 0.86fF
C20 n-leg_2/vpulldown n-leg_2/pd_ctrl 0.02fF
C21 p-leg_3/n_pu_ctrl p-leg_6/n_cal_ctrl[2] 0.25fF
C22 n-leg_3/pd_ctrl p-leg_6/n_cal_ctrl[2] 0.06fF
C23 p-leg_2/li_16_1957# n-leg_1/pd_ctrl 0.54fF
C24 p-leg_0/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.42fF
C25 p-leg_6/n_cal_ctrl[1] VDD 8.22fF
C26 p-leg_6/li_16_1957# p-leg_6/n_pu_ctrl 0.30fF
C27 pd_cal_ctrl[0] n-leg_1/pd_ctrl 0.11fF
C28 extr_sky130_fd_sc_hd__clkinv_4_4/Y VDD 0.15fF
C29 n-leg_0/vpulldown pd_cal_ctrl[0] 0.16fF
C30 p-leg_6/n_cal_ctrl[3] p-leg_6/li_16_1957# 0.17fF
C31 p-leg_6/n_cal_ctrl[2] VDD 8.10fF
C32 extr_sky130_fd_sc_hd__clkinv_4_7/Y p-leg_4/li_16_1957# 0.04fF
C33 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# p-leg_2/li_16_1957# 0.06fF
C34 extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47# p-leg_1/n_pu_ctrl 0.06fF
C35 pd_cal_ctrl[0] p-leg_4/li_16_1957# 0.66fF
C36 n-leg_1/vpulldown DQ 0.38fF
C37 p-leg_6/n_cal_ctrl[0] p-leg_0/n_pu_ctrl 0.58fF
C38 n-leg_1/vpulldown pd_cal_ctrl[2] 0.26fF
C39 pu_ctrl[5] extr_sky130_fd_sc_hd__clkbuf_16_5/X 0.03fF
C40 pd_cal_ctrl[3] n-leg_4/pd_ctrl 0.08fF
C41 extr_sky130_fd_sc_hd__clkinv_4_5/Y extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.03fF
C42 pd_cal_ctrl[0] n-leg_5/pd_ctrl 0.11fF
C43 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# n-leg_1/pd_ctrl 0.03fF
C44 VDD extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.13fF
C45 p-leg_2/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.38fF
C46 pd_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] 1.29fF
C47 DQ p-leg_1/n_pu_ctrl 0.71fF
C48 pu_cal_ctrl[2] p-leg_6/n_cal_ctrl[3] 0.03fF
C49 pd_cal_ctrl[3] p-leg_3/li_16_1957# 0.21fF
C50 p-leg_2/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.41fF
C51 extr_sky130_fd_sc_hd__clkbuf_16_6/X p-leg_6/li_16_1957# 0.04fF
C52 p-leg_2/n_pu_ctrl p-leg_6/n_cal_ctrl[1] 0.35fF
C53 pd_cal_ctrl[0] p-leg_6/n_cal_ctrl[2] 0.45fF
C54 pd_cal_ctrl[2] p-leg_1/n_pu_ctrl 0.25fF
C55 pd_ctrl[5] extr_sky130_fd_sc_hd__clkbuf_16_6/X 0.05fF
C56 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.05fF
C57 p-leg_6/n_cal_ctrl[2] p-leg_2/n_pu_ctrl 0.24fF
C58 n-leg_4/pd_ctrl VDD 0.06fF
C59 extr_sky130_fd_sc_hd__clkbuf_16_0/a_110_47# p-leg_0/n_pu_ctrl 0.06fF
C60 p-leg_3/n_pu_ctrl p-leg_3/li_16_1957# 0.30fF
C61 n-leg_1/pd_ctrl p-leg_6/n_cal_ctrl[2] 0.06fF
C62 p-leg_6/n_cal_ctrl[3] n-leg_0/pd_ctrl 0.21fF
C63 extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# pd_ctrl[2] 0.09fF
C64 pu_ctrl[3] VDD -0.03fF
C65 p-leg_4/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.38fF
C66 p-leg_3/li_16_1957# VDD 0.01fF
C67 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# p-leg_6/n_cal_ctrl[1] 0.21fF
C68 pu_cal_ctrl[3] VDD 0.39fF
C69 p-leg_1/extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C70 n-leg_1/vpulldown pd_cal_ctrl[1] 0.23fF
C71 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# p-leg_6/n_cal_ctrl[1] 0.21fF
C72 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.03fF
C73 p-leg_4/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.41fF
C74 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# p-leg_6/n_cal_ctrl[2] 0.17fF
C75 extr_sky130_fd_sc_hd__clkbuf_16_0/a_110_47# extr_sky130_fd_sc_hd__clkinv_16_2/A 0.26fF
C76 p-leg_5/n_pu_ctrl pd_cal_ctrl[3] 0.35fF
C77 extr_sky130_fd_sc_hd__clkbuf_16_5/X VDD 0.73fF
C78 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_4/Y 0.05fF
C79 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# p-leg_6/n_cal_ctrl[2] 0.17fF
C80 extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# n-leg_6/pd_ctrl 0.03fF
C81 DQ extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.03fF
C82 p-leg_6/n_cal_ctrl[2] n-leg_5/pd_ctrl 0.06fF
C83 pd_cal_ctrl[2] n-leg_6/vpulldown 0.08fF
C84 extr_sky130_fd_sc_hd__clkinv_4_4/Y p-leg_6/n_cal_ctrl[1] 0.09fF
C85 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_8/Y 0.17fF
C86 p-leg_1/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C87 pd_cal_ctrl[0] n-leg_4/pd_ctrl 0.11fF
C88 extr_sky130_fd_sc_hd__clkinv_4_6/Y extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.05fF
C89 pu_ctrl[0] extr_sky130_fd_sc_hd__clkinv_16_2/A 0.03fF
C90 p-leg_6/n_cal_ctrl[2] p-leg_6/n_cal_ctrl[1] 6.03fF
C91 pd_cal_ctrl[3] DQ 1.04fF
C92 p-leg_6/n_cal_ctrl[3] p-leg_5/li_16_1957# 0.38fF
C93 p-leg_6/n_cal_ctrl[3] p-leg_1/li_16_1957# 0.38fF
C94 p-leg_5/n_pu_ctrl VDD 0.76fF
C95 pd_cal_ctrl[0] p-leg_3/li_16_1957# 0.66fF
C96 extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47# extr_sky130_fd_sc_hd__clkinv_16_5/A 0.26fF
C97 p-leg_6/n_cal_ctrl[3] n-leg_2/pd_ctrl 0.21fF
C98 pd_cal_ctrl[3] pd_cal_ctrl[2] 17.76fF
C99 extr_sky130_fd_sc_hd__clkinv_16_8/A extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.26fF
C100 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# VDD 0.05fF
C101 DQ n-leg_3/pd_ctrl 0.11fF
C102 p-leg_3/n_pu_ctrl DQ 0.71fF
C103 pu_cal_ctrl[0] VDD 0.39fF
C104 p-leg_0/li_16_1957# DQ 0.28fF
C105 p-leg_6/n_cal_ctrl[0] pu_cal_ctrl[1] 0.08fF
C106 extr_sky130_fd_sc_hd__clkinv_4_9/Y extr_sky130_fd_sc_hd__clkinv_4_8/Y 0.28fF
C107 extr_sky130_fd_sc_hd__clkinv_4_9/Y pd_ctrl[4] 0.05fF
C108 p-leg_3/n_pu_ctrl pd_cal_ctrl[2] 0.25fF
C109 n-leg_3/pd_ctrl pd_cal_ctrl[2] 0.11fF
C110 DQ VDD 3.41fF
C111 p-leg_0/li_16_1957# pd_cal_ctrl[2] 0.29fF
C112 extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# VDD 0.05fF
C113 DQ extr_sky130_fd_sc_hd__clkinv_16_5/A 0.03fF
C114 pd_cal_ctrl[2] VDD 6.93fF
C115 pd_cal_ctrl[1] n-leg_6/vpulldown 0.09fF
C116 extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47# p-leg_4/n_pu_ctrl 0.06fF
C117 n-leg_3/vpulldown pd_cal_ctrl[3] 0.22fF
C118 p-leg_5/n_pu_ctrl pd_cal_ctrl[0] 0.86fF
C119 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# p-leg_3/li_16_1957# 0.06fF
C120 extr_sky130_fd_sc_hd__clkinv_4_13/Y pd_ctrl[6] 0.05fF
C121 p-leg_6/n_cal_ctrl[2] n-leg_4/pd_ctrl 0.06fF
C122 pd_cal_ctrl[3] pd_cal_ctrl[1] 7.04fF
C123 n-leg_3/vpulldown n-leg_3/pd_ctrl 0.02fF
C124 pu_cal_ctrl[3] p-leg_6/n_cal_ctrl[1] 0.02fF
C125 p-leg_3/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.38fF
C126 p-leg_2/li_16_1957# DQ 0.39fF
C127 p-leg_6/n_cal_ctrl[0] p-leg_1/n_pu_ctrl 0.58fF
C128 p-leg_3/li_16_1957# extr_sky130_fd_sc_hd__clkinv_4_4/Y 0.08fF
C129 pd_cal_ctrl[0] DQ 2.51fF
C130 extr_sky130_fd_sc_hd__clkinv_4_5/Y VDD 0.13fF
C131 p-leg_3/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.41fF
C132 pu_cal_ctrl[3] p-leg_6/n_cal_ctrl[2] 0.08fF
C133 pu_cal_ctrl[2] pu_cal_ctrl[1] 0.13fF
C134 p-leg_3/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C135 n-leg_3/pd_ctrl pd_cal_ctrl[1] 0.11fF
C136 DQ p-leg_2/n_pu_ctrl 0.71fF
C137 p-leg_2/li_16_1957# pd_cal_ctrl[2] 0.29fF
C138 p-leg_3/extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C139 p-leg_0/li_16_1957# pd_cal_ctrl[1] 0.25fF
C140 pd_cal_ctrl[0] pd_cal_ctrl[2] 7.42fF
C141 extr_sky130_fd_sc_hd__clkinv_4_1/Y VDD 0.13fF
C142 n-leg_1/pd_ctrl DQ 0.11fF
C143 pd_cal_ctrl[1] VDD 7.47fF
C144 pd_cal_ctrl[2] p-leg_2/n_pu_ctrl 0.25fF
C145 extr_sky130_fd_sc_hd__clkinv_4_1/Y extr_sky130_fd_sc_hd__clkinv_16_5/A 0.10fF
C146 n-leg_0/vpulldown DQ 0.38fF
C147 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.17fF
C148 n-leg_1/pd_ctrl pd_cal_ctrl[2] 0.11fF
C149 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# VDD 0.05fF
C150 n-leg_0/vpulldown pd_cal_ctrl[2] 0.26fF
C151 DQ p-leg_4/li_16_1957# 0.39fF
C152 p-leg_5/n_pu_ctrl p-leg_6/n_cal_ctrl[1] 0.35fF
C153 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# n-leg_5/pd_ctrl 0.03fF
C154 p-leg_6/li_16_1957# extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.08fF
C155 p-leg_6/n_cal_ctrl[3] p-leg_4/n_pu_ctrl 0.25fF
C156 p-leg_5/li_16_1957# extr_sky130_fd_sc_hd__clkinv_4_8/Y 0.08fF
C157 p-leg_5/n_pu_ctrl p-leg_6/n_cal_ctrl[2] 0.24fF
C158 pd_ctrl[5] extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.01fF
C159 pd_cal_ctrl[2] p-leg_4/li_16_1957# 0.29fF
C160 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# p-leg_6/n_cal_ctrl[1] 0.21fF
C161 pu_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] 0.03fF
C162 pd_cal_ctrl[0] n-leg_3/vpulldown 0.16fF
C163 DQ n-leg_5/pd_ctrl 0.11fF
C164 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# p-leg_6/n_cal_ctrl[2] 0.17fF
C165 extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47# pd_ctrl[4] 0.09fF
C166 p-leg_2/li_16_1957# pd_cal_ctrl[1] 0.25fF
C167 DQ p-leg_6/n_cal_ctrl[1] 1.10fF
C168 p-leg_6/n_cal_ctrl[1] extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.21fF
C169 pd_ctrl[5] extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.09fF
C170 pd_cal_ctrl[2] n-leg_5/pd_ctrl 0.11fF
C171 pd_cal_ctrl[0] pd_cal_ctrl[1] 18.62fF
C172 p-leg_6/n_cal_ctrl[0] pd_cal_ctrl[3] 1.63fF
C173 DQ p-leg_6/n_cal_ctrl[2] 1.35fF
C174 p-leg_6/n_cal_ctrl[3] p-leg_0/n_pu_ctrl 0.25fF
C175 pd_cal_ctrl[2] p-leg_6/n_cal_ctrl[1] 1.62fF
C176 p-leg_6/n_cal_ctrl[2] extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.17fF
C177 p-leg_2/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C178 pd_ctrl[3] extr_sky130_fd_sc_hd__clkinv_4_6/Y 0.01fF
C179 extr_sky130_fd_sc_hd__clkbuf_16_6/X p-leg_6/n_pu_ctrl 1.37fF
C180 n-leg_1/pd_ctrl pd_cal_ctrl[1] 0.11fF
C181 pd_cal_ctrl[2] p-leg_6/n_cal_ctrl[2] 0.45fF
C182 extr_sky130_fd_sc_hd__clkinv_4_0/Y VDD 0.15fF
C183 pd_cal_ctrl[3] p-leg_6/li_16_1957# 0.21fF
C184 n-leg_3/vpulldown p-leg_4/li_16_1957# 0.60fF
C185 p-leg_6/n_cal_ctrl[0] p-leg_3/n_pu_ctrl 0.58fF
C186 p-leg_6/n_cal_ctrl[0] n-leg_3/pd_ctrl 0.21fF
C187 n-leg_0/vpulldown pd_cal_ctrl[1] 0.23fF
C188 p-leg_6/n_cal_ctrl[0] p-leg_0/li_16_1957# 0.39fF
C189 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.01fF
C190 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C191 extr_sky130_fd_sc_hd__clkinv_4_13/Y VDD 0.13fF
C192 p-leg_6/n_cal_ctrl[0] VDD 8.20fF
C193 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_3/Y 0.19fF
C194 p-leg_4/li_16_1957# pd_cal_ctrl[1] 0.25fF
C195 extr_sky130_fd_sc_hd__clkinv_4_5/Y extr_sky130_fd_sc_hd__clkinv_4_4/Y 0.28fF
C196 p-leg_6/li_16_1957# VDD 0.01fF
C197 pd_cal_ctrl[1] n-leg_5/pd_ctrl 0.11fF
C198 pd_cal_ctrl[3] n-leg_4/vpulldown 0.22fF
C199 extr_sky130_fd_sc_hd__clkinv_4_6/Y VDD 0.15fF
C200 p-leg_6/n_cal_ctrl[1] pd_cal_ctrl[1] 1.29fF
C201 extr_sky130_fd_sc_hd__clkinv_16_2/A p-leg_0/n_pu_ctrl 1.37fF
C202 DQ n-leg_4/pd_ctrl 0.11fF
C203 p-leg_1/n_pu_ctrl p-leg_1/li_16_1957# 0.30fF
C204 p-leg_5/n_pu_ctrl extr_sky130_fd_sc_hd__clkbuf_16_5/X 1.37fF
C205 n-leg_4/pd_ctrl extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.03fF
C206 extr_sky130_fd_sc_hd__clkinv_4_9/Y VDD 0.13fF
C207 p-leg_6/n_cal_ctrl[2] pd_cal_ctrl[1] 0.45fF
C208 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# p-leg_6/n_cal_ctrl[1] 0.21fF
C209 pd_cal_ctrl[2] n-leg_4/pd_ctrl 0.11fF
C210 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_7/Y 0.19fF
C211 p-leg_6/n_cal_ctrl[0] p-leg_2/li_16_1957# 0.38fF
C212 p-leg_6/n_cal_ctrl[3] extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.17fF
C213 p-leg_3/li_16_1957# DQ 0.39fF
C214 p-leg_6/n_cal_ctrl[0] pd_cal_ctrl[0] 1.30fF
C215 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# p-leg_6/n_cal_ctrl[2] 0.17fF
C216 pd_cal_ctrl[3] n-leg_0/pd_ctrl 0.08fF
C217 extr_sky130_fd_sc_hd__clkinv_4_4/Y pd_ctrl[2] 0.01fF
C218 p-leg_6/n_cal_ctrl[0] p-leg_2/n_pu_ctrl 0.58fF
C219 DQ extr_sky130_fd_sc_hd__clkbuf_16_5/X 0.03fF
C220 p-leg_3/li_16_1957# pd_cal_ctrl[2] 0.29fF
C221 pu_cal_ctrl[2] VDD 0.39fF
C222 extr_sky130_fd_sc_hd__clkinv_16_9/A extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.31fF
C223 pd_cal_ctrl[0] p-leg_6/li_16_1957# 0.66fF
C224 p-leg_6/n_cal_ctrl[0] n-leg_1/pd_ctrl 0.21fF
C225 extr_sky130_fd_sc_hd__clkinv_4_6/Y extr_sky130_fd_sc_hd__clkinv_4_7/Y 0.28fF
C226 n-leg_6/pd_ctrl n-leg_6/vpulldown 0.02fF
C227 extr_sky130_fd_sc_hd__clkbuf_8_6/A extr_sky130_fd_sc_hd__clkinv_4_13/Y 0.28fF
C228 extr_sky130_fd_sc_hd__clkinv_4_2/Y VDD 0.15fF
C229 extr_sky130_fd_sc_hd__clkinv_4_3/Y extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.28fF
C230 pd_ctrl[1] extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C231 p-leg_6/n_cal_ctrl[0] p-leg_4/li_16_1957# 0.38fF
C232 pd_cal_ctrl[3] n-leg_2/vpulldown 0.22fF
C233 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# p-leg_6/n_cal_ctrl[0] 0.03fF
C234 n-leg_0/pd_ctrl VDD 0.06fF
C235 p-leg_5/n_pu_ctrl DQ 0.71fF
C236 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# p-leg_6/n_cal_ctrl[0] 0.03fF
C237 extr_sky130_fd_sc_hd__clkinv_4_5/Y p-leg_3/li_16_1957# 0.04fF
C238 extr_sky130_fd_sc_hd__clkinv_16_8/A VDD 0.73fF
C239 extr_sky130_fd_sc_hd__clkinv_4_0/Y p-leg_6/n_cal_ctrl[1] 0.09fF
C240 extr_sky130_fd_sc_hd__clkinv_4_3/Y extr_sky130_fd_sc_hd__clkinv_16_8/A 0.10fF
C241 extr_sky130_fd_sc_hd__clkinv_16_5/A pd_ctrl[0] 0.05fF
C242 n-leg_5/vpulldown pd_cal_ctrl[3] 0.22fF
C243 n-leg_4/pd_ctrl pd_cal_ctrl[1] 0.11fF
C244 extr_sky130_fd_sc_hd__clkinv_16_8/A pd_ctrl[1] 0.05fF
C245 p-leg_5/n_pu_ctrl pd_cal_ctrl[2] 0.25fF
C246 pd_cal_ctrl[3] p-leg_5/li_16_1957# 0.21fF
C247 pd_cal_ctrl[0] n-leg_4/vpulldown 0.16fF
C248 p-leg_6/n_cal_ctrl[0] n-leg_5/pd_ctrl 0.21fF
C249 pd_cal_ctrl[3] p-leg_1/li_16_1957# 0.21fF
C250 extr_sky130_fd_sc_hd__clkinv_4_6/Y p-leg_4/li_16_1957# 0.08fF
C251 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] 7.02fF
C252 pd_cal_ctrl[3] n-leg_2/pd_ctrl 0.08fF
C253 p-leg_3/li_16_1957# pd_cal_ctrl[1] 0.25fF
C254 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_4/Y 0.17fF
C255 n-leg_6/pd_ctrl VDD 0.06fF
C256 p-leg_6/li_16_1957# n-leg_5/pd_ctrl 0.54fF
C257 p-leg_2/li_16_1957# extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.08fF
C258 p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[2] 1.30fF
C259 DQ pd_cal_ctrl[2] 0.86fF
C260 p-leg_6/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.07fF
C261 p-leg_5/li_16_1957# VDD 0.01fF
C262 p-leg_6/extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C263 extr_sky130_fd_sc_hd__clkinv_4_6/Y p-leg_6/n_cal_ctrl[1] 0.09fF
C264 extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47# extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.26fF
C265 pd_cal_ctrl[0] n-leg_0/pd_ctrl 0.11fF
C266 pd_ctrl[3] extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.11fF
C267 p-leg_1/li_16_1957# VDD 0.01fF
C268 p-leg_6/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.20fF
C269 p-leg_2/li_16_1957# extr_sky130_fd_sc_hd__clkinv_16_8/A 0.04fF
C270 VDD n-leg_2/pd_ctrl 0.06fF
C271 extr_sky130_fd_sc_hd__clkinv_16_5/A p-leg_1/li_16_1957# 0.04fF
C272 extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_1/Y 0.03fF
C273 p-leg_6/n_cal_ctrl[3] p-leg_1/n_pu_ctrl 0.25fF
C274 extr_sky130_fd_sc_hd__clkinv_16_8/A p-leg_2/n_pu_ctrl 1.37fF
C275 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.19fF
C276 p-leg_5/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C277 n-leg_0/vpulldown n-leg_0/pd_ctrl 0.02fF
C278 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.05fF
C279 pd_cal_ctrl[0] n-leg_2/vpulldown 0.16fF
C280 n-leg_3/vpulldown DQ 0.38fF
C281 p-leg_6/li_16_1957# extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.04fF
C282 pu_cal_ctrl[2] p-leg_6/n_cal_ctrl[1] 0.08fF
C283 pd_ctrl[5] extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.05fF
C284 n-leg_5/vpulldown pd_cal_ctrl[0] 0.16fF
C285 n-leg_3/vpulldown pd_cal_ctrl[2] 0.26fF
C286 pd_cal_ctrl[0] p-leg_5/li_16_1957# 0.66fF
C287 p-leg_6/n_cal_ctrl[0] n-leg_4/pd_ctrl 0.21fF
C288 pu_cal_ctrl[2] p-leg_6/n_cal_ctrl[2] 0.19fF
C289 DQ pd_cal_ctrl[1] 2.08fF
C290 pd_cal_ctrl[0] p-leg_1/li_16_1957# 0.66fF
C291 p-leg_6/n_cal_ctrl[1] extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.09fF
C292 pu_ctrl[1] extr_sky130_fd_sc_hd__clkinv_16_5/A 0.03fF
C293 extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47# p-leg_6/n_pu_ctrl 0.06fF
C294 pd_cal_ctrl[0] n-leg_2/pd_ctrl 0.11fF
C295 extr_sky130_fd_sc_hd__clkinv_16_8/A pu_ctrl[2] 0.03fF
C296 extr_sky130_fd_sc_hd__clkinv_4_8/Y pd_ctrl[4] 0.01fF
C297 pd_cal_ctrl[2] pd_cal_ctrl[1] 17.82fF
C298 p-leg_6/n_cal_ctrl[0] p-leg_3/li_16_1957# 0.38fF
C299 n-leg_0/vpulldown p-leg_1/li_16_1957# 0.60fF
C300 n-leg_0/pd_ctrl p-leg_6/n_cal_ctrl[2] 0.06fF
C301 p-leg_4/n_pu_ctrl extr_sky130_fd_sc_hd__clkbuf_16_4/X 1.37fF
C302 extr_sky130_fd_sc_hd__clkinv_16_9/A p-leg_3/n_pu_ctrl 1.37fF
C303 pd_cal_ctrl[3] p-leg_6/n_pu_ctrl 0.35fF
C304 p-leg_6/n_cal_ctrl[3] pd_cal_ctrl[3] 0.45fF
C305 pd_cal_ctrl[3] p-leg_4/n_pu_ctrl 0.35fF
C306 extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_7/Y 0.03fF
C307 extr_sky130_fd_sc_hd__clkinv_16_9/A VDD 0.75fF
C308 n-leg_5/vpulldown n-leg_5/pd_ctrl 0.02fF
C309 n-leg_4/pd_ctrl n-leg_4/vpulldown 0.02fF
C310 n-leg_3/vpulldown pd_cal_ctrl[1] 0.23fF
C311 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# n-leg_2/pd_ctrl 0.03fF
C312 p-leg_6/n_cal_ctrl[0] p-leg_5/n_pu_ctrl 0.58fF
C313 extr_sky130_fd_sc_hd__clkinv_4_9/Y extr_sky130_fd_sc_hd__clkbuf_16_5/X 0.10fF
C314 p-leg_6/n_cal_ctrl[3] p-leg_3/n_pu_ctrl 0.25fF
C315 p-leg_6/n_cal_ctrl[3] n-leg_3/pd_ctrl 0.21fF
C316 p-leg_5/li_16_1957# p-leg_6/n_cal_ctrl[1] 0.38fF
C317 p-leg_0/li_16_1957# p-leg_6/n_cal_ctrl[3] 0.39fF
C318 extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47# extr_sky130_fd_sc_hd__clkbuf_16_6/X 0.31fF
C319 p-leg_6/n_pu_ctrl VDD 0.76fF
C320 p-leg_6/n_cal_ctrl[1] p-leg_1/li_16_1957# 0.38fF
C321 extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# VDD 0.05fF
C322 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# p-leg_6/n_cal_ctrl[0] 0.03fF
C323 pu_cal_ctrl[0] p-leg_6/n_cal_ctrl[0] 0.20fF
C324 p-leg_5/li_16_1957# p-leg_6/n_cal_ctrl[2] 0.41fF
C325 extr_sky130_fd_sc_hd__clkinv_4_1/Y extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# 0.01fF
C326 pd_cal_ctrl[3] p-leg_0/n_pu_ctrl 0.35fF
C327 pu_cal_ctrl[3] pu_cal_ctrl[2] 0.13fF
C328 p-leg_6/n_cal_ctrl[3] VDD 7.52fF
C329 p-leg_4/n_pu_ctrl VDD 0.76fF
C330 extr_sky130_fd_sc_hd__clkinv_4_5/Y pd_ctrl[2] 0.05fF
C331 p-leg_6/n_cal_ctrl[2] p-leg_1/li_16_1957# 0.41fF
C332 p-leg_6/n_cal_ctrl[2] n-leg_2/pd_ctrl 0.06fF
C333 p-leg_6/n_cal_ctrl[0] DQ 1.68fF
C334 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.03fF
C335 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# p-leg_6/li_16_1957# 0.06fF
C336 p-leg_0/li_16_1957# p-leg_0/n_pu_ctrl 0.30fF
C337 p-leg_6/n_cal_ctrl[0] pd_cal_ctrl[2] 1.63fF
C338 p-leg_6/li_16_1957# DQ 0.39fF
C339 p-leg_0/n_pu_ctrl VDD 0.76fF
C340 p-leg_6/li_16_1957# pd_cal_ctrl[2] 0.29fF
C341 pd_cal_ctrl[0] p-leg_6/n_pu_ctrl 0.86fF
C342 p-leg_2/li_16_1957# p-leg_6/n_cal_ctrl[3] 0.38fF
C343 p-leg_0/li_16_1957# extr_sky130_fd_sc_hd__clkinv_16_2/A 0.04fF
C344 extr_sky130_fd_sc_hd__clkinv_4_9/Y extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.01fF
C345 pd_cal_ctrl[0] p-leg_6/n_cal_ctrl[3] 0.45fF
C346 extr_sky130_fd_sc_hd__clkbuf_16_6/X VDD 0.77fF
C347 pd_cal_ctrl[0] p-leg_4/n_pu_ctrl 0.86fF
C348 extr_sky130_fd_sc_hd__clkinv_4_3/Y extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.03fF
C349 extr_sky130_fd_sc_hd__clkinv_4_1/Y extr_sky130_fd_sc_hd__clkinv_4_0/Y 0.28fF
C350 pd_ctrl[1] extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.09fF
C351 extr_sky130_fd_sc_hd__clkinv_16_2/A VDD 0.73fF
C352 n-leg_2/vpulldown p-leg_3/li_16_1957# 0.60fF
C353 p-leg_6/n_cal_ctrl[3] p-leg_2/n_pu_ctrl 0.25fF
C354 p-leg_5/li_16_1957# n-leg_4/pd_ctrl 0.54fF
C355 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_5/Y 0.19fF
C356 extr_sky130_fd_sc_hd__clkbuf_16_6/X pu_ctrl[6] 0.04fF
C357 DQ n-leg_4/vpulldown 0.38fF
C358 p-leg_6/n_cal_ctrl[3] n-leg_1/pd_ctrl 0.21fF
C359 extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47# pd_ctrl[0] 0.11fF
C360 extr_sky130_fd_sc_hd__clkinv_4_1/Y p-leg_6/n_cal_ctrl[0] 0.19fF
C361 extr_sky130_fd_sc_hd__clkinv_4_0/Y extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# 0.05fF
C362 extr_sky130_fd_sc_hd__clkbuf_8_6/A extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# 0.05fF
C363 pd_cal_ctrl[2] n-leg_4/vpulldown 0.26fF
C364 p-leg_6/n_cal_ctrl[0] pd_cal_ctrl[1] 1.30fF
C365 pd_cal_ctrl[0] p-leg_0/n_pu_ctrl 0.86fF
C366 p-leg_6/n_cal_ctrl[3] p-leg_4/li_16_1957# 0.38fF
C367 p-leg_3/li_16_1957# n-leg_2/pd_ctrl 0.54fF
C368 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# p-leg_6/n_cal_ctrl[3] 0.17fF
C369 p-leg_5/li_16_1957# extr_sky130_fd_sc_hd__clkbuf_16_5/X 0.04fF
C370 p-leg_4/li_16_1957# p-leg_4/n_pu_ctrl 0.30fF
C371 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# 0.03fF
C372 n-leg_3/pd_ctrl extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.03fF
C373 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# p-leg_6/n_cal_ctrl[3] 0.17fF
C374 p-leg_6/li_16_1957# pd_cal_ctrl[1] 0.25fF
C375 DQ n-leg_0/pd_ctrl 0.11fF
C376 extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47# extr_sky130_fd_sc_hd__clkbuf_16_5/X 0.26fF
C377 p-leg_6/n_cal_ctrl[3] n-leg_5/pd_ctrl 0.21fF
C378 VDD extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.05fF
C379 extr_sky130_fd_sc_hd__clkinv_16_8/A DQ 0.03fF
C380 extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47# p-leg_2/n_pu_ctrl 0.06fF
C381 pd_cal_ctrl[2] n-leg_0/pd_ctrl 0.11fF
C382 p-leg_6/n_cal_ctrl[3] p-leg_6/n_cal_ctrl[1] 1.69fF
C383 p-leg_4/n_pu_ctrl p-leg_6/n_cal_ctrl[1] 0.35fF
C384 p-leg_5/n_pu_ctrl p-leg_5/li_16_1957# 0.30fF
C385 p-leg_6/n_cal_ctrl[3] p-leg_6/n_cal_ctrl[2] 5.56fF
C386 p-leg_4/n_pu_ctrl p-leg_6/n_cal_ctrl[2] 0.24fF
C387 extr_sky130_fd_sc_hd__clkinv_4_8/Y VDD 0.15fF
C388 n-leg_2/vpulldown DQ 0.38fF
C389 extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47# p-leg_5/n_pu_ctrl 0.06fF
C390 n-leg_4/vpulldown pd_cal_ctrl[1] 0.23fF
C391 p-leg_3/n_pu_ctrl extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.06fF
C392 n-leg_5/vpulldown DQ 0.38fF
C393 n-leg_2/vpulldown pd_cal_ctrl[2] 0.26fF
C394 p-leg_5/li_16_1957# DQ 0.39fF
C395 p-leg_6/n_cal_ctrl[1] p-leg_0/n_pu_ctrl 0.35fF
C396 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_0/Y 0.17fF
C397 p-leg_5/li_16_1957# extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.06fF
C398 DQ p-leg_1/li_16_1957# 0.39fF
C399 extr_sky130_fd_sc_hd__clkinv_4_7/Y extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.01fF
C400 extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VDD -0.06fF
C401 n-leg_1/vpulldown pd_cal_ctrl[3] 0.22fF
C402 n-leg_5/vpulldown pd_cal_ctrl[2] 0.26fF
C403 DQ n-leg_2/pd_ctrl 0.11fF
C404 p-leg_6/n_cal_ctrl[2] p-leg_0/n_pu_ctrl 0.24fF
C405 p-leg_5/li_16_1957# pd_cal_ctrl[2] 0.29fF
C406 pu_cal_ctrl[1] VDD 0.39fF
C407 pd_cal_ctrl[2] p-leg_1/li_16_1957# 0.29fF
C408 extr_sky130_fd_sc_hd__clkinv_4_1/Y pd_ctrl[0] 0.05fF
C409 p-leg_0/extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C410 pd_cal_ctrl[2] n-leg_2/pd_ctrl 0.11fF
C411 n-leg_0/pd_ctrl pd_cal_ctrl[1] 0.11fF
C412 extr_sky130_fd_sc_hd__clkinv_16_9/A pu_ctrl[3] 0.04fF
C413 extr_sky130_fd_sc_hd__clkinv_16_9/A p-leg_3/li_16_1957# 0.04fF
C414 pd_cal_ctrl[3] p-leg_1/n_pu_ctrl 0.35fF
C415 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# n-leg_0/pd_ctrl 0.03fF
C416 p-leg_6/n_cal_ctrl[0] p-leg_6/li_16_1957# 0.07fF
C417 p-leg_6/n_cal_ctrl[3] n-leg_4/pd_ctrl 0.21fF
C418 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_6/Y 0.17fF
C419 p-leg_4/li_16_1957# extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.06fF
C420 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_9/Y 0.19fF
C421 n-leg_2/vpulldown pd_cal_ctrl[1] 0.29fF
C422 p-leg_6/n_cal_ctrl[3] p-leg_3/li_16_1957# 0.38fF
C423 pu_cal_ctrl[3] p-leg_6/n_cal_ctrl[3] 0.19fF
C424 extr_sky130_fd_sc_hd__clkbuf_16_6/X extr_sky130_fd_sc_hd__clkinv_4_11/Y 0.10fF
C425 n-leg_5/vpulldown pd_cal_ctrl[1] 0.29fF
C426 extr_sky130_fd_sc_hd__clkinv_4_1/Y p-leg_1/li_16_1957# 0.04fF
C427 p-leg_1/n_pu_ctrl VDD 0.77fF
C428 p-leg_5/li_16_1957# pd_cal_ctrl[1] 0.25fF
C429 p-leg_6/n_cal_ctrl[1] extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.21fF
C430 p-leg_1/li_16_1957# pd_cal_ctrl[1] 0.25fF
C431 extr_sky130_fd_sc_hd__clkinv_16_5/A p-leg_1/n_pu_ctrl 1.38fF
C432 p-leg_6/n_cal_ctrl[0] pu_cal_ctrl[2] 0.02fF
C433 pd_cal_ctrl[1] n-leg_2/pd_ctrl 0.11fF
C434 pd_ctrl[3] extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.05fF
C435 p-leg_6/n_cal_ctrl[2] extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# 0.17fF
C436 p-leg_2/li_16_1957# n-leg_1/vpulldown 0.60fF
C437 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# p-leg_1/li_16_1957# 0.06fF
C438 n-leg_1/vpulldown pd_cal_ctrl[0] 0.16fF
C439 pd_cal_ctrl[3] n-leg_6/vpulldown 0.03fF
C440 extr_sky130_fd_sc_hd__clkinv_4_0/Y pd_ctrl[0] 0.01fF
C441 p-leg_6/n_cal_ctrl[1] extr_sky130_fd_sc_hd__clkinv_4_8/Y 0.09fF
C442 VDD extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.15fF
C443 p-leg_6/n_cal_ctrl[0] extr_sky130_fd_sc_hd__clkinv_4_2/Y 0.17fF
C444 extr_sky130_fd_sc_hd__clkinv_16_9/A DQ 0.03fF
C445 p-leg_5/n_pu_ctrl p-leg_6/n_cal_ctrl[3] 0.25fF
C446 pu_ctrl[4] extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.03fF
C447 n-leg_1/vpulldown n-leg_1/pd_ctrl 0.02fF
C448 p-leg_6/n_cal_ctrl[0] n-leg_0/pd_ctrl 0.21fF
C449 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# p-leg_6/n_cal_ctrl[3] 0.17fF
C450 pd_cal_ctrl[0] p-leg_1/n_pu_ctrl 0.86fF
C451 DQ p-leg_6/n_pu_ctrl 0.71fF
C452 p-leg_6/n_cal_ctrl[3] DQ 1.23fF
C453 DQ p-leg_4/n_pu_ctrl 0.71fF
C454 p-leg_6/n_cal_ctrl[3] extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# 0.17fF
C455 VDD extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.73fF
C456 p-leg_6/n_cal_ctrl[1] pu_cal_ctrl[1] 0.19fF
C457 pd_cal_ctrl[3] p-leg_3/n_pu_ctrl 0.35fF
C458 pd_cal_ctrl[2] p-leg_6/n_pu_ctrl 0.25fF
C459 pd_cal_ctrl[3] n-leg_3/pd_ctrl 0.08fF
C460 p-leg_0/li_16_1957# pd_cal_ctrl[3] 0.21fF
C461 p-leg_6/n_cal_ctrl[3] pd_cal_ctrl[2] 0.45fF
C462 p-leg_6/n_cal_ctrl[2] pu_cal_ctrl[1] 0.03fF
C463 pd_cal_ctrl[2] p-leg_4/n_pu_ctrl 0.25fF
C464 extr_sky130_fd_sc_hd__clkbuf_8_6/A pd_ctrl[6] 0.01fF
C465 extr_sky130_fd_sc_hd__clkinv_4_0/Y p-leg_1/li_16_1957# 0.08fF
C466 pd_cal_ctrl[3] VDD 7.04fF
C467 extr_sky130_fd_sc_hd__clkinv_4_5/Y extr_sky130_fd_sc_hd__clkinv_16_9/A 0.10fF
C468 p-leg_6/n_cal_ctrl[0] p-leg_5/li_16_1957# 0.38fF
C469 DQ p-leg_0/n_pu_ctrl 0.71fF
C470 p-leg_6/n_cal_ctrl[0] p-leg_1/li_16_1957# 0.38fF
C471 n-leg_3/pd_ctrl VDD 0.06fF
C472 p-leg_3/n_pu_ctrl VDD 0.76fF
C473 p-leg_6/n_cal_ctrl[0] n-leg_2/pd_ctrl 0.21fF
C474 p-leg_0/li_16_1957# VDD 0.01fF
C475 n-leg_5/vpulldown p-leg_6/li_16_1957# 0.60fF
C476 pd_cal_ctrl[2] p-leg_0/n_pu_ctrl 0.24fF
C477 pd_cal_ctrl[0] n-leg_6/vpulldown 0.06fF
C478 extr_sky130_fd_sc_hd__clkinv_4_7/Y extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.10fF
C479 pd_ctrl[3] extr_sky130_fd_sc_hd__clkinv_4_7/Y 0.05fF
C480 extr_sky130_fd_sc_hd__clkbuf_16_6/X DQ 0.03fF
C481 extr_sky130_fd_sc_hd__clkinv_4_3/Y VDD 0.13fF
C482 p-leg_1/n_pu_ctrl p-leg_6/n_cal_ctrl[1] 0.35fF
C483 extr_sky130_fd_sc_hd__clkinv_4_3/Y pd_ctrl[1] 0.05fF
C484 DQ extr_sky130_fd_sc_hd__clkinv_16_2/A 0.03fF
C485 extr_sky130_fd_sc_hd__clkinv_16_5/A VDD 0.73fF
C486 p-leg_6/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C487 p-leg_5/li_16_1957# extr_sky130_fd_sc_hd__clkinv_4_9/Y 0.04fF
C488 p-leg_2/li_16_1957# pd_cal_ctrl[3] 0.21fF
C489 p-leg_6/n_cal_ctrl[2] p-leg_1/n_pu_ctrl 0.24fF
C490 pd_cal_ctrl[0] pd_cal_ctrl[3] 5.32fF
C491 extr_sky130_fd_sc_hd__clkinv_16_9/A pd_ctrl[2] 0.05fF
C492 p-leg_6/n_cal_ctrl[3] pd_cal_ctrl[1] 0.45fF
C493 p-leg_4/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C494 extr_sky130_fd_sc_hd__clkbuf_16_5/X pd_ctrl[4] 0.05fF
C495 pd_cal_ctrl[3] p-leg_2/n_pu_ctrl 0.35fF
C496 extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47# extr_sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C497 p-leg_4/extr_sky130_fd_sc_hd__fill_8_9/VPWR VDD 0.55fF
C498 p-leg_6/n_cal_ctrl[3] extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# 0.17fF
C499 p-leg_5/li_16_1957# n-leg_4/vpulldown 0.60fF
C500 p-leg_6/n_cal_ctrl[1] extr_sky130_fd_sc_hd__clkbuf_8_5/A 0.09fF
C501 pd_cal_ctrl[0] p-leg_3/n_pu_ctrl 0.86fF
C502 n-leg_1/pd_ctrl pd_cal_ctrl[3] 0.08fF
C503 pd_cal_ctrl[0] n-leg_3/pd_ctrl 0.11fF
C504 p-leg_0/li_16_1957# pd_cal_ctrl[0] 0.66fF
C505 p-leg_4/li_16_1957# extr_sky130_fd_sc_hd__clkbuf_16_4/X 0.04fF
C506 n-leg_0/vpulldown pd_cal_ctrl[3] 0.22fF
C507 extr_sky130_fd_sc_hd__clkinv_4_7/Y VDD 0.13fF
C508 p-leg_2/li_16_1957# VDD 0.01fF
C509 extr_sky130_fd_sc_hd__clkinv_4_3/Y p-leg_2/li_16_1957# 0.04fF
C510 pd_cal_ctrl[0] VDD 6.93fF
C511 p-leg_0/n_pu_ctrl pd_cal_ctrl[1] 0.38fF
C512 pd_cal_ctrl[3] p-leg_4/li_16_1957# 0.21fF
C513 p-leg_2/n_pu_ctrl VDD 0.76fF
C514 n-leg_1/pd_ctrl VDD 0.06fF
C515 n-leg_0/pd_ctrl p-leg_1/li_16_1957# 0.54fF
C516 pd_cal_ctrl[3] n-leg_5/pd_ctrl 0.08fF
C517 n-leg_3/pd_ctrl p-leg_4/li_16_1957# 0.54fF
C518 n-leg_0/pd_ctrl GND 8.25fF
C519 extr_sky130_fd_sc_hd__clkinv_4_0/Y GND 0.23fF
C520 extr_sky130_fd_sc_hd__clkbuf_8_0/a_110_47# GND 0.94fF
C521 p-leg_2/li_16_1957# GND -6.69fF
C522 p-leg_2/n_pu_ctrl GND 3.53fF
C523 pu_cal_ctrl[3] GND 0.07fF
C524 pu_cal_ctrl[2] GND 0.06fF
C525 p-leg_1/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND 0.16fF
C526 p-leg_1/li_16_1957# GND -6.69fF
C527 p-leg_1/n_pu_ctrl GND 3.49fF
C528 p-leg_0/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND 0.16fF
C529 p-leg_0/li_16_1957# GND -6.69fF
C530 p-leg_0/n_pu_ctrl GND 3.53fF
C531 pu_cal_ctrl[1] GND 0.07fF
C532 pu_cal_ctrl[0] GND 0.06fF
C533 pu_ctrl[6] GND 0.61fF
C534 extr_sky130_fd_sc_hd__clkbuf_16_6/a_110_47# GND 1.83fF
C535 pu_ctrl[5] GND 0.59fF
C536 extr_sky130_fd_sc_hd__clkbuf_16_5/a_110_47# GND 1.83fF
C537 pu_ctrl[4] GND 0.59fF
C538 extr_sky130_fd_sc_hd__clkbuf_16_4/a_110_47# GND 1.83fF
C539 pu_ctrl[3] GND 0.64fF
C540 extr_sky130_fd_sc_hd__clkbuf_16_3/a_110_47# GND 1.83fF
C541 pu_ctrl[2] GND 0.59fF
C542 extr_sky130_fd_sc_hd__clkbuf_16_2/a_110_47# GND 1.83fF
C543 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND 5.92fF
C544 pu_ctrl[1] GND 0.59fF
C545 extr_sky130_fd_sc_hd__clkbuf_16_1/a_110_47# GND 1.83fF
C546 pu_ctrl[0] GND 0.60fF
C547 extr_sky130_fd_sc_hd__clkbuf_16_0/a_110_47# GND 1.84fF
C548 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND 6.13fF
C549 pd_ctrl[4] GND 0.67fF
C550 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND 5.89fF
C551 extr_sky130_fd_sc_hd__clkinv_4_9/Y GND 0.68fF
C552 pd_ctrl[3] GND 0.65fF
C553 extr_sky130_fd_sc_hd__clkinv_16_9/A GND 5.96fF
C554 extr_sky130_fd_sc_hd__clkinv_4_7/Y GND 0.60fF
C555 pd_ctrl[2] GND 0.71fF
C556 extr_sky130_fd_sc_hd__clkinv_4_5/Y GND 0.81fF
C557 extr_sky130_fd_sc_hd__clkinv_16_8/A GND 6.13fF
C558 pd_ctrl[1] GND 0.67fF
C559 extr_sky130_fd_sc_hd__clkinv_4_3/Y GND 0.67fF
C560 extr_sky130_fd_sc_hd__clkinv_4_1/Y GND 0.60fF
C561 pd_ctrl[0] GND 0.65fF
C562 extr_sky130_fd_sc_hd__clkinv_16_5/A GND 5.88fF
C563 n-leg_6/vpulldown GND 11.94fF
C564 pd_cal_ctrl[1] GND 18.00fF
C565 pd_cal_ctrl[3] GND 16.32fF
C566 pd_cal_ctrl[0] GND 30.53fF
C567 pd_cal_ctrl[2] GND 14.44fF
C568 pd_ctrl[6] GND 0.71fF
C569 n-leg_6/pd_ctrl GND 8.39fF
C570 extr_sky130_fd_sc_hd__clkbuf_8_6/A GND 0.38fF
C571 extr_sky130_fd_sc_hd__clkbuf_8_6/a_110_47# GND 0.94fF
C572 n-leg_5/vpulldown GND 11.94fF
C573 extr_sky130_fd_sc_hd__clkinv_4_13/Y GND 0.81fF
C574 n-leg_5/pd_ctrl GND 8.39fF
C575 extr_sky130_fd_sc_hd__clkbuf_8_5/A GND 0.38fF
C576 extr_sky130_fd_sc_hd__clkbuf_8_5/a_110_47# GND 0.94fF
C577 n-leg_4/vpulldown GND 11.94fF
C578 pd_ctrl[5] GND 0.71fF
C579 n-leg_4/pd_ctrl GND 8.31fF
C580 extr_sky130_fd_sc_hd__clkinv_4_8/Y GND 0.27fF
C581 extr_sky130_fd_sc_hd__clkbuf_8_4/a_110_47# GND 0.94fF
C582 extr_sky130_fd_sc_hd__clkinv_16_2/A GND 5.97fF
C583 p-leg_6/n_cal_ctrl[1] GND -4.41fF
C584 VDD GND 371.65fF
C585 p-leg_6/n_cal_ctrl[3] GND 10.78fF
C586 p-leg_6/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND 0.16fF
C587 p-leg_6/n_cal_ctrl[2] GND -3.89fF
C588 DQ GND -22.45fF
C589 p-leg_6/li_16_1957# GND -6.69fF
C590 p-leg_6/n_cal_ctrl[0] GND -1.36fF
C591 p-leg_6/n_pu_ctrl GND 3.54fF
C592 n-leg_3/vpulldown GND 11.94fF
C593 extr_sky130_fd_sc_hd__clkinv_4_11/Y GND 0.81fF
C594 n-leg_3/pd_ctrl GND 8.25fF
C595 extr_sky130_fd_sc_hd__clkinv_4_6/Y GND 0.23fF
C596 extr_sky130_fd_sc_hd__clkbuf_8_3/a_110_47# GND 0.94fF
C597 p-leg_5/li_16_1957# GND -6.69fF
C598 p-leg_5/n_pu_ctrl GND 3.53fF
C599 n-leg_2/vpulldown GND 11.94fF
C600 n-leg_2/pd_ctrl GND 8.39fF
C601 extr_sky130_fd_sc_hd__clkinv_4_4/Y GND 0.38fF
C602 extr_sky130_fd_sc_hd__clkbuf_8_2/a_110_47# GND 0.94fF
C603 p-leg_4/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND 0.16fF
C604 p-leg_4/li_16_1957# GND -6.69fF
C605 p-leg_4/n_pu_ctrl GND 3.42fF
C606 n-leg_1/vpulldown GND 11.94fF
C607 n-leg_1/pd_ctrl GND 8.30fF
C608 extr_sky130_fd_sc_hd__clkinv_4_2/Y GND 0.26fF
C609 extr_sky130_fd_sc_hd__clkbuf_8_1/a_110_47# GND 0.94fF
C610 p-leg_3/extr_sky130_fd_sc_hd__fill_8_9/VPWR GND 0.16fF
C611 p-leg_3/li_16_1957# GND -6.69fF
C612 p-leg_3/n_pu_ctrl GND 3.52fF
C613 n-leg_0/vpulldown GND 11.94fF
.ends

