magic
tech sky130A
magscale 1 2
timestamp 1644036613
<< viali >>
rect 5 222 50 267
rect 281 214 315 248
rect 1477 222 1522 267
rect 1753 214 1787 248
rect 2949 222 2994 267
rect 3225 214 3259 248
rect 4421 222 4466 267
rect 4697 214 4731 248
rect 5893 222 5938 267
rect 6169 214 6203 248
rect 7365 222 7410 267
rect 7641 214 7675 248
rect 8837 222 8882 267
rect 9113 214 9147 248
rect 10585 214 10619 248
rect 1370 101 1411 142
rect 2842 101 2883 142
rect 4314 101 4355 142
rect 5786 101 5827 142
rect 7258 101 7299 142
rect 8730 101 8771 142
rect 10202 101 10243 142
rect 11674 101 11715 142
<< metal1 >>
rect -1 267 56 279
rect 1471 267 1528 279
rect 2943 267 3000 279
rect 4415 267 4472 279
rect 5887 267 5944 279
rect 7359 267 7416 279
rect 8831 267 8888 279
rect -50 222 5 267
rect 50 248 1477 267
rect 50 222 281 248
rect -1 210 56 222
rect 275 214 281 222
rect 315 222 1477 248
rect 1522 248 2949 267
rect 1522 222 1753 248
rect 315 214 321 222
rect 275 202 321 214
rect 1471 210 1528 222
rect 1747 214 1753 222
rect 1787 222 2949 248
rect 2994 248 4421 267
rect 2994 222 3225 248
rect 1787 214 1793 222
rect 1747 202 1793 214
rect 2943 210 3000 222
rect 3219 214 3225 222
rect 3259 222 4421 248
rect 4466 248 5893 267
rect 4466 222 4697 248
rect 3259 214 3265 222
rect 3219 202 3265 214
rect 4415 210 4472 222
rect 4691 214 4697 222
rect 4731 222 5893 248
rect 5938 248 7365 267
rect 5938 222 6169 248
rect 4731 214 4737 222
rect 4691 202 4737 214
rect 5887 210 5944 222
rect 6163 214 6169 222
rect 6203 222 7365 248
rect 7410 248 8837 267
rect 7410 222 7641 248
rect 6203 214 6209 222
rect 6163 202 6209 214
rect 7359 210 7416 222
rect 7635 214 7641 222
rect 7675 222 8837 248
rect 8882 248 11802 267
rect 8882 222 9113 248
rect 7675 214 7681 222
rect 7635 202 7681 214
rect 8831 210 8888 222
rect 9107 214 9113 222
rect 9147 222 10585 248
rect 9147 214 9153 222
rect 9107 202 9153 214
rect 10579 214 10585 222
rect 10619 222 11802 248
rect 10619 214 10625 222
rect 10579 202 10625 214
rect 277 142 318 202
rect -12 101 318 142
rect 1364 148 1458 154
rect 1364 142 1406 148
rect 1749 142 1790 202
rect 1364 101 1370 142
rect 1458 101 1790 142
rect 2836 148 2930 154
rect 2836 142 2878 148
rect 3221 142 3262 202
rect 2836 101 2842 142
rect 2930 101 3262 142
rect 4308 148 4402 154
rect 4308 142 4350 148
rect 4693 142 4734 202
rect 4308 101 4314 142
rect 4402 101 4734 142
rect 5780 148 5874 154
rect 5780 142 5822 148
rect 6165 142 6206 202
rect 5780 101 5786 142
rect 5874 101 6206 142
rect 7252 148 7346 154
rect 7252 142 7294 148
rect 7637 142 7678 202
rect 7252 101 7258 142
rect 7346 101 7678 142
rect 8724 148 8818 154
rect 8724 142 8766 148
rect 9109 142 9150 202
rect 8724 101 8730 142
rect 8818 101 9150 142
rect 10196 148 10290 154
rect 10196 142 10238 148
rect 10581 142 10622 202
rect 10196 101 10202 142
rect 10290 101 10622 142
rect 11668 148 11762 154
rect 11668 142 11710 148
rect 11668 101 11674 142
rect 11762 101 11802 142
rect 1364 96 1406 101
rect 1364 90 1458 96
rect 2836 96 2878 101
rect 2836 90 2930 96
rect 4308 96 4350 101
rect 4308 90 4402 96
rect 5780 96 5822 101
rect 5780 90 5874 96
rect 7252 96 7294 101
rect 7252 90 7346 96
rect 8724 96 8766 101
rect 8724 90 8818 96
rect 10196 96 10238 101
rect 10196 90 10290 96
rect 11668 96 11710 101
rect 11668 90 11762 96
rect 1364 89 1417 90
rect 2836 89 2889 90
rect 4308 89 4361 90
rect 5780 89 5833 90
rect 7252 89 7305 90
rect 8724 89 8777 90
rect 10196 89 10249 90
rect 11668 89 11721 90
<< via1 >>
rect 1406 142 1458 148
rect 1406 101 1411 142
rect 1411 101 1458 142
rect 2878 142 2930 148
rect 2878 101 2883 142
rect 2883 101 2930 142
rect 4350 142 4402 148
rect 4350 101 4355 142
rect 4355 101 4402 142
rect 5822 142 5874 148
rect 5822 101 5827 142
rect 5827 101 5874 142
rect 7294 142 7346 148
rect 7294 101 7299 142
rect 7299 101 7346 142
rect 8766 142 8818 148
rect 8766 101 8771 142
rect 8771 101 8818 142
rect 10238 142 10290 148
rect 10238 101 10243 142
rect 10243 101 10290 142
rect 11710 142 11762 148
rect 11710 101 11715 142
rect 11715 101 11762 142
rect 1406 96 1458 101
rect 2878 96 2930 101
rect 4350 96 4402 101
rect 5822 96 5874 101
rect 7294 96 7346 101
rect 8766 96 8818 101
rect 10238 96 10290 101
rect 11710 96 11762 101
<< metal2 >>
rect 1412 148 1452 604
rect 2884 148 2924 604
rect 4356 148 4396 604
rect 5828 148 5868 604
rect 7300 148 7340 604
rect 8772 148 8812 604
rect 10244 148 10284 604
rect 11716 148 11756 604
rect 1400 96 1406 148
rect 1458 96 1464 148
rect 2872 96 2878 148
rect 2930 96 2936 148
rect 4344 96 4350 148
rect 4402 96 4408 148
rect 5816 96 5822 148
rect 5874 96 5880 148
rect 7288 96 7294 148
rect 7346 96 7352 148
rect 8760 96 8766 148
rect 8818 96 8824 148
rect 10232 96 10238 148
rect 10290 96 10296 148
rect 11704 96 11710 148
rect 11762 96 11768 148
rect 1412 -36 1452 96
rect 2884 -36 2924 96
rect 4356 -36 4396 96
rect 5828 -36 5868 96
rect 7300 -36 7340 96
rect 8772 -36 8812 96
rect 10244 -36 10284 96
rect 11716 -36 11756 96
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7 ~/cad/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1643856600
transform 1 0 10292 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1643856600
transform 1 0 8820 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1643856600
transform 1 0 7348 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1643856600
transform 1 0 5876 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1643856600
transform 1 0 4404 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1643856600
transform 1 0 2932 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1643856600
transform 1 0 1460 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1643856600
transform 1 0 -12 0 1 12
box -38 -48 1510 592
<< end >>
