magic
tech sky130A
magscale 1 2
timestamp 1646981735
<< poly >>
rect 2301 221 2331 289
<< locali >>
rect 3910 2004 3957 2031
rect 2481 872 2637 913
rect 4228 861 4340 895
rect 5976 861 6088 895
rect 7724 861 7836 895
rect 9472 861 9584 895
rect 11220 861 11332 895
rect 12968 861 13080 895
rect 14716 861 14828 895
rect 4309 699 4388 767
rect 4456 699 4527 767
rect 2206 308 2343 361
rect 200 188 388 294
rect 476 188 665 294
rect 752 188 943 294
rect 1134 233 1172 307
rect 2206 291 2273 308
rect 1376 250 1497 284
rect 1652 253 1774 287
rect 1928 257 2053 291
rect 3938 262 4032 311
rect 5686 262 5780 311
rect 7434 262 7528 311
rect 9182 262 9276 311
rect 10930 262 11024 311
rect 12678 262 12772 311
rect 14426 262 14520 311
rect 2273 231 2343 238
rect 3940 247 3987 262
rect 3940 203 3941 247
rect 3985 203 3987 247
rect 3940 202 3987 203
rect 5688 247 5735 262
rect 5688 203 5689 247
rect 5733 203 5735 247
rect 5688 202 5735 203
rect 7436 247 7483 262
rect 7436 203 7437 247
rect 7481 203 7483 247
rect 7436 202 7483 203
rect 9184 247 9231 262
rect 9184 203 9185 247
rect 9229 203 9231 247
rect 9184 202 9231 203
rect 10932 247 10979 262
rect 10932 203 10933 247
rect 10977 203 10979 247
rect 10932 202 10979 203
rect 12680 247 12727 262
rect 12680 203 12681 247
rect 12725 203 12727 247
rect 12680 202 12727 203
rect 14428 247 14475 262
rect 14428 203 14429 247
rect 14473 203 14475 247
rect 14428 202 14475 203
rect 532 -222 722 -116
rect 809 -222 998 -116
<< viali >>
rect 3731 1978 3787 2034
rect 3910 1957 3957 2004
rect 4119 1963 4154 1998
rect 3288 1549 3322 1583
rect 4313 1549 4347 1583
rect 6057 1549 6091 1583
rect 9468 1549 9502 1583
rect 3207 1413 3241 1447
rect 4400 1413 4434 1447
rect 6148 1413 6182 1447
rect 3115 1324 3155 1364
rect 4120 1342 4160 1382
rect 5878 1342 5918 1382
rect 7792 1345 7826 1379
rect 7878 1342 7918 1382
rect 7982 1342 8022 1382
rect 9370 1345 9404 1379
rect 9651 1342 9691 1382
rect 11296 1342 11336 1382
rect 11384 1345 11418 1379
rect 11478 1342 11518 1382
rect 13042 1342 13082 1382
rect 13138 1345 13172 1379
rect 13229 1342 13269 1382
rect 14886 1342 14926 1382
rect 15038 1345 15072 1379
rect 15165 1342 15205 1382
rect 3491 1261 3525 1295
rect 4688 1267 4722 1301
rect 6436 1267 6470 1301
rect 8160 1229 8218 1287
rect 9932 1267 9966 1301
rect 11656 1229 11714 1287
rect 13404 1229 13462 1287
rect 15155 1217 15189 1251
rect 2279 867 2337 925
rect 2749 888 2805 944
rect 3488 876 3528 916
rect 4037 882 4077 922
rect 4685 860 4725 900
rect 5785 882 5825 922
rect 6433 860 6473 900
rect 7533 882 7573 922
rect 9281 882 9321 922
rect 8166 824 8212 870
rect 9929 860 9969 900
rect 11029 882 11069 922
rect 12777 882 12817 922
rect 11662 824 11708 870
rect 14525 882 14565 922
rect 13410 824 13456 870
rect 15152 822 15192 862
rect 4388 699 4456 767
rect 6135 705 6191 761
rect 7922 705 7978 761
rect 9641 705 9697 761
rect 11372 705 11428 761
rect 13127 705 13183 761
rect 14884 705 14940 761
rect 66 254 113 301
rect 1060 234 1099 273
rect 2273 238 2343 308
rect 4032 262 4081 311
rect 5780 262 5829 311
rect 7528 262 7577 311
rect 9276 262 9325 311
rect 11024 262 11073 311
rect 12772 262 12821 311
rect 14520 262 14569 311
rect 2529 197 2585 253
rect 3941 203 3985 247
rect 4277 197 4333 253
rect 5689 203 5733 247
rect 6025 197 6081 253
rect 7437 203 7481 247
rect 7773 197 7829 253
rect 9185 203 9229 247
rect 9521 197 9577 253
rect 10933 203 10977 247
rect 11269 197 11325 253
rect 12681 203 12725 247
rect 13017 197 13073 253
rect 14429 203 14473 247
rect 344 -222 403 -116
rect 1118 -221 1158 -181
<< metal1 >>
rect 3719 1972 3725 2040
rect 3793 1972 3799 2040
rect 3898 2004 3969 2010
rect 3898 1957 3910 2004
rect 3957 1998 4166 2004
rect 3957 1963 4119 1998
rect 4154 1963 4166 1998
rect 3957 1957 4166 1963
rect 3898 1951 3969 1957
rect 3276 1583 3334 1589
rect 4108 1583 4114 1592
rect 47 1552 3288 1583
rect 47 1549 3081 1552
rect 3189 1549 3288 1552
rect 3322 1549 4114 1583
rect 3276 1543 3334 1549
rect 4108 1540 4114 1549
rect 4166 1540 4172 1592
rect 4301 1583 4359 1592
rect 4301 1549 4313 1583
rect 4347 1549 4359 1583
rect 3103 1515 3109 1524
rect 47 1481 3109 1515
rect 3103 1472 3109 1481
rect 3161 1515 3167 1524
rect 4301 1515 4359 1549
rect 4485 1540 4491 1592
rect 4543 1583 4549 1592
rect 6045 1583 6103 1589
rect 7970 1583 7976 1592
rect 4543 1552 6057 1583
rect 4543 1549 5838 1552
rect 5958 1549 6057 1552
rect 6091 1552 7976 1583
rect 6091 1549 7844 1552
rect 7952 1549 7976 1552
rect 4543 1540 4549 1549
rect 6045 1543 6103 1549
rect 7970 1540 7976 1549
rect 8028 1583 8034 1592
rect 9462 1583 9508 1589
rect 11466 1583 11472 1592
rect 8028 1549 9468 1583
rect 9502 1552 11472 1583
rect 9502 1549 9617 1552
rect 9725 1549 11256 1552
rect 11376 1549 11472 1552
rect 8028 1540 8034 1549
rect 9462 1543 9508 1549
rect 11466 1540 11472 1549
rect 11524 1583 11530 1592
rect 13030 1583 13036 1592
rect 11524 1549 13036 1583
rect 11524 1540 11530 1549
rect 13030 1540 13036 1549
rect 13088 1583 13094 1592
rect 15153 1583 15159 1592
rect 13088 1552 15159 1583
rect 13088 1549 13195 1552
rect 13303 1549 14852 1552
rect 14960 1549 15159 1552
rect 13088 1540 13094 1549
rect 15153 1540 15159 1549
rect 15211 1583 15217 1592
rect 15211 1549 15227 1583
rect 15211 1540 15217 1549
rect 5866 1515 5872 1524
rect 3161 1512 4080 1515
rect 4200 1512 4457 1515
rect 4577 1512 5872 1515
rect 3161 1481 5872 1512
rect 3161 1472 3167 1481
rect 5866 1472 5872 1481
rect 5924 1515 5930 1524
rect 7866 1515 7872 1524
rect 5924 1481 7872 1515
rect 5924 1472 5930 1481
rect 7866 1472 7872 1481
rect 7924 1515 7930 1524
rect 9639 1515 9645 1524
rect 7924 1512 7942 1515
rect 8062 1512 9645 1515
rect 7924 1481 9645 1512
rect 7924 1472 7930 1481
rect 9639 1472 9645 1481
rect 9697 1515 9703 1524
rect 11284 1515 11290 1524
rect 9697 1481 11290 1515
rect 9697 1472 9703 1481
rect 11284 1472 11290 1481
rect 11342 1515 11348 1524
rect 13217 1515 13223 1524
rect 11342 1512 11444 1515
rect 11564 1512 13008 1515
rect 13116 1512 13223 1515
rect 11342 1481 13223 1512
rect 11342 1472 11348 1481
rect 13217 1472 13223 1481
rect 13275 1515 13281 1524
rect 14874 1515 14880 1524
rect 13275 1481 14880 1515
rect 13275 1472 13281 1481
rect 14874 1472 14880 1481
rect 14932 1515 14938 1524
rect 14932 1512 15131 1515
rect 14932 1481 15227 1512
rect 14932 1472 14938 1481
rect 3195 1447 3253 1453
rect 4388 1447 4446 1453
rect 6136 1447 6194 1453
rect 47 1444 3081 1447
rect 3189 1444 3207 1447
rect 47 1413 3207 1444
rect 3241 1416 4400 1447
rect 3241 1413 4080 1416
rect 4200 1413 4400 1416
rect 4434 1444 5838 1447
rect 5958 1444 6148 1447
rect 4434 1416 6148 1444
rect 4434 1413 5838 1416
rect 5958 1413 6148 1416
rect 6182 1444 7844 1447
rect 7964 1444 9617 1447
rect 9725 1444 11256 1447
rect 11376 1444 13195 1447
rect 13303 1444 14852 1447
rect 14960 1444 15227 1447
rect 6182 1416 15227 1444
rect 6182 1413 7838 1416
rect 8062 1413 9611 1416
rect 9731 1413 11256 1416
rect 11376 1413 11438 1416
rect 11558 1413 13002 1416
rect 13110 1413 13201 1416
rect 13309 1413 14846 1416
rect 14966 1413 15125 1416
rect 3195 1407 3253 1413
rect 4388 1407 4446 1413
rect 6136 1407 6194 1413
rect 3103 1318 3109 1370
rect 3161 1318 3167 1370
rect 4108 1333 4114 1388
rect 4166 1376 4172 1388
rect 4485 1376 4491 1385
rect 4166 1342 4491 1376
rect 4166 1333 4172 1342
rect 4485 1333 4491 1342
rect 4543 1333 4549 1385
rect 5866 1336 5872 1388
rect 5924 1336 5930 1388
rect 7786 1379 7832 1413
rect 7786 1345 7792 1379
rect 7826 1345 7832 1379
rect 7786 1333 7832 1345
rect 7866 1336 7872 1388
rect 7924 1336 7930 1388
rect 7970 1336 7976 1388
rect 8028 1336 8034 1388
rect 9364 1379 9410 1413
rect 9364 1345 9370 1379
rect 9404 1345 9410 1379
rect 9364 1333 9410 1345
rect 9639 1336 9645 1388
rect 9697 1336 9703 1388
rect 11284 1336 11290 1388
rect 11342 1336 11348 1388
rect 11378 1379 11424 1413
rect 11378 1345 11384 1379
rect 11418 1345 11424 1379
rect 11378 1333 11424 1345
rect 11466 1336 11472 1388
rect 11524 1336 11530 1388
rect 13030 1336 13036 1388
rect 13088 1336 13094 1388
rect 13132 1379 13178 1413
rect 13132 1345 13138 1379
rect 13172 1345 13178 1379
rect 13132 1333 13178 1345
rect 13217 1336 13223 1388
rect 13275 1336 13281 1388
rect 14874 1336 14880 1388
rect 14932 1336 14938 1388
rect 15032 1379 15078 1413
rect 15032 1345 15038 1379
rect 15072 1345 15078 1379
rect 15032 1333 15078 1345
rect 15153 1336 15159 1388
rect 15211 1336 15217 1388
rect 4679 1310 4731 1316
rect 3482 1304 3534 1310
rect 4679 1252 4731 1258
rect 6427 1310 6479 1316
rect 9923 1310 9975 1316
rect 6427 1252 6479 1258
rect 8148 1293 8230 1299
rect 3482 1246 3534 1252
rect 8148 1223 8154 1293
rect 8224 1223 8230 1293
rect 9923 1252 9975 1258
rect 11644 1293 11726 1299
rect 8148 1217 8230 1223
rect 11644 1223 11650 1293
rect 11720 1223 11726 1293
rect 11644 1217 11726 1223
rect 13392 1293 13474 1299
rect 13392 1223 13398 1293
rect 13468 1223 13474 1293
rect 13392 1217 13474 1223
rect 15146 1260 15198 1266
rect 15146 1202 15198 1208
rect 2743 944 2811 956
rect 2267 861 2273 931
rect 2343 861 2349 931
rect 2743 888 2749 944
rect 2805 888 2811 944
rect 2743 767 2811 888
rect 3476 870 3482 922
rect 3534 870 3540 922
rect 4025 876 4031 928
rect 4083 876 4089 928
rect 4673 854 4679 906
rect 4731 854 4737 906
rect 5773 876 5779 928
rect 5831 876 5837 928
rect 6421 854 6427 906
rect 6479 854 6485 906
rect 7521 876 7527 928
rect 7579 876 7585 928
rect 9269 876 9275 928
rect 9327 876 9333 928
rect 8154 818 8160 876
rect 8218 818 8224 876
rect 9917 854 9923 906
rect 9975 854 9981 906
rect 11017 876 11023 928
rect 11075 876 11081 928
rect 12765 876 12771 928
rect 12823 876 12829 928
rect 14513 876 14519 928
rect 14571 876 14577 928
rect 11650 818 11656 876
rect 11714 818 11720 876
rect 13398 818 13404 876
rect 13462 818 13468 876
rect 15140 816 15146 868
rect 15198 816 15204 868
rect 3725 767 3793 773
rect 4382 767 4462 779
rect 2743 699 3725 767
rect 3793 699 4388 767
rect 4456 761 15019 767
rect 4456 705 6135 761
rect 6191 705 7922 761
rect 7978 705 9641 761
rect 9697 705 11372 761
rect 11428 705 13127 761
rect 13183 705 14884 761
rect 14940 705 15019 761
rect 4456 699 15019 705
rect 3725 693 3793 699
rect 4382 687 4462 699
rect 2261 314 2355 320
rect 54 248 60 307
rect 119 248 125 307
rect 1048 273 1112 279
rect 1048 234 1060 273
rect 1099 234 1112 273
rect 1048 228 1112 234
rect 1106 227 1112 228
rect 1164 227 1170 279
rect 2261 232 2267 314
rect 2349 232 2355 314
rect 4026 317 4087 323
rect 5774 317 5835 323
rect 7522 317 7583 323
rect 9270 317 9331 323
rect 11018 317 11079 323
rect 12766 317 12827 323
rect 14514 317 14575 323
rect 2261 226 2355 232
rect 2523 253 2591 265
rect 4026 262 4032 265
rect 4081 262 4087 265
rect 2523 197 2529 253
rect 2585 247 3997 253
rect 4026 250 4087 262
rect 4271 253 4339 265
rect 5774 262 5780 265
rect 5829 262 5835 265
rect 2585 203 3941 247
rect 3985 203 3997 247
rect 2585 197 3997 203
rect 4271 197 4277 253
rect 4333 247 5745 253
rect 5774 250 5835 262
rect 6019 253 6087 265
rect 7522 262 7528 265
rect 7577 262 7583 265
rect 4333 203 5689 247
rect 5733 203 5745 247
rect 4333 197 5745 203
rect 6019 197 6025 253
rect 6081 247 7493 253
rect 7522 250 7583 262
rect 7767 253 7835 265
rect 9270 262 9276 265
rect 9325 262 9331 265
rect 6081 203 7437 247
rect 7481 203 7493 247
rect 6081 197 7493 203
rect 7767 197 7773 253
rect 7829 247 9241 253
rect 9270 250 9331 262
rect 9515 253 9583 265
rect 11018 262 11024 265
rect 11073 262 11079 265
rect 7829 203 9185 247
rect 9229 203 9241 247
rect 7829 197 9241 203
rect 9515 197 9521 253
rect 9577 247 10989 253
rect 11018 250 11079 262
rect 11263 253 11331 265
rect 12766 262 12772 265
rect 12821 262 12827 265
rect 9577 203 10933 247
rect 10977 203 10989 247
rect 9577 197 10989 203
rect 11263 197 11269 253
rect 11325 247 12737 253
rect 12766 250 12827 262
rect 13011 253 13079 265
rect 14514 262 14520 265
rect 14569 262 14575 265
rect 11325 203 12681 247
rect 12725 203 12737 247
rect 11325 197 12737 203
rect 13011 197 13017 253
rect 13073 247 14485 253
rect 14514 250 14575 262
rect 13073 203 14429 247
rect 14473 203 14485 247
rect 13073 197 14485 203
rect 2523 185 2591 197
rect 4271 185 4339 197
rect 6019 185 6087 197
rect 7767 185 7835 197
rect 9515 185 9583 197
rect 11263 185 11331 197
rect 13011 185 13079 197
rect 338 -116 409 -104
rect 338 -139 344 -116
rect 54 -198 60 -139
rect 119 -198 344 -139
rect 338 -222 344 -198
rect 403 -222 409 -116
rect 338 -234 409 -222
rect 1106 -227 1112 -175
rect 1164 -227 1170 -175
<< via1 >>
rect 3725 2034 3793 2040
rect 3725 1978 3731 2034
rect 3731 1978 3787 2034
rect 3787 1978 3793 2034
rect 3725 1972 3793 1978
rect 4114 1540 4166 1592
rect 3109 1472 3161 1524
rect 4491 1540 4543 1592
rect 7976 1540 8028 1592
rect 11472 1540 11524 1592
rect 13036 1540 13088 1592
rect 15159 1540 15211 1592
rect 5872 1472 5924 1524
rect 7872 1472 7924 1524
rect 9645 1472 9697 1524
rect 11290 1472 11342 1524
rect 13223 1472 13275 1524
rect 14880 1472 14932 1524
rect 3109 1364 3161 1370
rect 3109 1324 3115 1364
rect 3115 1324 3155 1364
rect 3155 1324 3161 1364
rect 3109 1318 3161 1324
rect 4114 1382 4166 1388
rect 4114 1342 4120 1382
rect 4120 1342 4160 1382
rect 4160 1342 4166 1382
rect 4114 1333 4166 1342
rect 4491 1333 4543 1385
rect 5872 1382 5924 1388
rect 5872 1342 5878 1382
rect 5878 1342 5918 1382
rect 5918 1342 5924 1382
rect 5872 1336 5924 1342
rect 7872 1382 7924 1388
rect 7872 1342 7878 1382
rect 7878 1342 7918 1382
rect 7918 1342 7924 1382
rect 7872 1336 7924 1342
rect 7976 1382 8028 1388
rect 7976 1342 7982 1382
rect 7982 1342 8022 1382
rect 8022 1342 8028 1382
rect 7976 1336 8028 1342
rect 9645 1382 9697 1388
rect 9645 1342 9651 1382
rect 9651 1342 9691 1382
rect 9691 1342 9697 1382
rect 9645 1336 9697 1342
rect 11290 1382 11342 1388
rect 11290 1342 11296 1382
rect 11296 1342 11336 1382
rect 11336 1342 11342 1382
rect 11290 1336 11342 1342
rect 11472 1382 11524 1388
rect 11472 1342 11478 1382
rect 11478 1342 11518 1382
rect 11518 1342 11524 1382
rect 11472 1336 11524 1342
rect 13036 1382 13088 1388
rect 13036 1342 13042 1382
rect 13042 1342 13082 1382
rect 13082 1342 13088 1382
rect 13036 1336 13088 1342
rect 13223 1382 13275 1388
rect 13223 1342 13229 1382
rect 13229 1342 13269 1382
rect 13269 1342 13275 1382
rect 13223 1336 13275 1342
rect 14880 1382 14932 1388
rect 14880 1342 14886 1382
rect 14886 1342 14926 1382
rect 14926 1342 14932 1382
rect 14880 1336 14932 1342
rect 15159 1382 15211 1388
rect 15159 1342 15165 1382
rect 15165 1342 15205 1382
rect 15205 1342 15211 1382
rect 15159 1336 15211 1342
rect 3482 1295 3534 1304
rect 3482 1261 3491 1295
rect 3491 1261 3525 1295
rect 3525 1261 3534 1295
rect 3482 1252 3534 1261
rect 4679 1301 4731 1310
rect 4679 1267 4688 1301
rect 4688 1267 4722 1301
rect 4722 1267 4731 1301
rect 4679 1258 4731 1267
rect 6427 1301 6479 1310
rect 6427 1267 6436 1301
rect 6436 1267 6470 1301
rect 6470 1267 6479 1301
rect 9923 1301 9975 1310
rect 6427 1258 6479 1267
rect 8154 1287 8224 1293
rect 8154 1229 8160 1287
rect 8160 1229 8218 1287
rect 8218 1229 8224 1287
rect 8154 1223 8224 1229
rect 9923 1267 9932 1301
rect 9932 1267 9966 1301
rect 9966 1267 9975 1301
rect 9923 1258 9975 1267
rect 11650 1287 11720 1293
rect 11650 1229 11656 1287
rect 11656 1229 11714 1287
rect 11714 1229 11720 1287
rect 11650 1223 11720 1229
rect 13398 1287 13468 1293
rect 13398 1229 13404 1287
rect 13404 1229 13462 1287
rect 13462 1229 13468 1287
rect 13398 1223 13468 1229
rect 15146 1251 15198 1260
rect 15146 1217 15155 1251
rect 15155 1217 15189 1251
rect 15189 1217 15198 1251
rect 15146 1208 15198 1217
rect 2273 925 2343 931
rect 2273 867 2279 925
rect 2279 867 2337 925
rect 2337 867 2343 925
rect 2273 861 2343 867
rect 3482 916 3534 922
rect 3482 876 3488 916
rect 3488 876 3528 916
rect 3528 876 3534 916
rect 3482 870 3534 876
rect 4031 922 4083 928
rect 4031 882 4037 922
rect 4037 882 4077 922
rect 4077 882 4083 922
rect 4031 876 4083 882
rect 4679 900 4731 906
rect 4679 860 4685 900
rect 4685 860 4725 900
rect 4725 860 4731 900
rect 4679 854 4731 860
rect 5779 922 5831 928
rect 5779 882 5785 922
rect 5785 882 5825 922
rect 5825 882 5831 922
rect 5779 876 5831 882
rect 6427 900 6479 906
rect 6427 860 6433 900
rect 6433 860 6473 900
rect 6473 860 6479 900
rect 6427 854 6479 860
rect 7527 922 7579 928
rect 7527 882 7533 922
rect 7533 882 7573 922
rect 7573 882 7579 922
rect 7527 876 7579 882
rect 9275 922 9327 928
rect 9275 882 9281 922
rect 9281 882 9321 922
rect 9321 882 9327 922
rect 9275 876 9327 882
rect 8160 870 8218 876
rect 8160 824 8166 870
rect 8166 824 8212 870
rect 8212 824 8218 870
rect 8160 818 8218 824
rect 9923 900 9975 906
rect 9923 860 9929 900
rect 9929 860 9969 900
rect 9969 860 9975 900
rect 9923 854 9975 860
rect 11023 922 11075 928
rect 11023 882 11029 922
rect 11029 882 11069 922
rect 11069 882 11075 922
rect 11023 876 11075 882
rect 12771 922 12823 928
rect 12771 882 12777 922
rect 12777 882 12817 922
rect 12817 882 12823 922
rect 12771 876 12823 882
rect 14519 922 14571 928
rect 14519 882 14525 922
rect 14525 882 14565 922
rect 14565 882 14571 922
rect 14519 876 14571 882
rect 11656 870 11714 876
rect 11656 824 11662 870
rect 11662 824 11708 870
rect 11708 824 11714 870
rect 11656 818 11714 824
rect 13404 870 13462 876
rect 13404 824 13410 870
rect 13410 824 13456 870
rect 13456 824 13462 870
rect 13404 818 13462 824
rect 15146 862 15198 868
rect 15146 822 15152 862
rect 15152 822 15192 862
rect 15192 822 15198 862
rect 15146 816 15198 822
rect 3725 699 3793 767
rect 60 301 119 307
rect 60 254 66 301
rect 66 254 113 301
rect 113 254 119 301
rect 60 248 119 254
rect 1112 227 1164 279
rect 2267 308 2349 314
rect 2267 238 2273 308
rect 2273 238 2343 308
rect 2343 238 2349 308
rect 2267 232 2349 238
rect 4026 311 4087 317
rect 4026 265 4032 311
rect 4032 265 4081 311
rect 4081 265 4087 311
rect 5774 311 5835 317
rect 5774 265 5780 311
rect 5780 265 5829 311
rect 5829 265 5835 311
rect 7522 311 7583 317
rect 7522 265 7528 311
rect 7528 265 7577 311
rect 7577 265 7583 311
rect 9270 311 9331 317
rect 9270 265 9276 311
rect 9276 265 9325 311
rect 9325 265 9331 311
rect 11018 311 11079 317
rect 11018 265 11024 311
rect 11024 265 11073 311
rect 11073 265 11079 311
rect 12766 311 12827 317
rect 12766 265 12772 311
rect 12772 265 12821 311
rect 12821 265 12827 311
rect 14514 311 14575 317
rect 14514 265 14520 311
rect 14520 265 14569 311
rect 14569 265 14575 311
rect 60 -198 119 -139
rect 1112 -181 1164 -175
rect 1112 -221 1118 -181
rect 1118 -221 1158 -181
rect 1158 -221 1164 -181
rect 1112 -227 1164 -221
<< metal2 >>
rect 3725 2040 3793 2046
rect 3103 1472 3109 1524
rect 3161 1472 3167 1524
rect 3118 1376 3152 1472
rect 3109 1370 3161 1376
rect 3109 1312 3161 1318
rect 3482 1304 3534 1310
rect 3482 1246 3534 1252
rect 2273 931 2343 937
rect 3491 928 3525 1246
rect 3482 922 3534 928
rect 3482 864 3534 870
rect 2273 320 2343 861
rect 3491 858 3525 864
rect 3725 767 3793 1972
rect 4114 1592 4166 1598
rect 4114 1534 4166 1540
rect 4491 1592 4543 1598
rect 4491 1534 4543 1540
rect 7976 1592 8028 1598
rect 11466 1540 11472 1592
rect 11524 1540 11530 1592
rect 13030 1540 13036 1592
rect 13088 1540 13094 1592
rect 15153 1540 15159 1592
rect 15211 1540 15217 1592
rect 7976 1534 8028 1540
rect 4123 1394 4157 1534
rect 4114 1388 4166 1394
rect 4500 1391 4534 1534
rect 5872 1524 5924 1530
rect 7866 1472 7872 1524
rect 7924 1472 7930 1524
rect 5872 1466 5924 1472
rect 5881 1394 5915 1466
rect 7881 1394 7915 1472
rect 7985 1394 8019 1534
rect 11290 1524 11342 1530
rect 9639 1472 9645 1524
rect 9697 1472 9703 1524
rect 9654 1394 9688 1472
rect 11290 1466 11342 1472
rect 11299 1394 11333 1466
rect 11481 1394 11515 1540
rect 13045 1394 13079 1540
rect 13217 1472 13223 1524
rect 13275 1472 13281 1524
rect 14874 1472 14880 1524
rect 14932 1472 14938 1524
rect 13232 1394 13266 1472
rect 14889 1394 14923 1472
rect 15168 1394 15202 1540
rect 4114 1327 4166 1333
rect 4491 1385 4543 1391
rect 4491 1327 4543 1333
rect 5872 1388 5924 1394
rect 5872 1330 5924 1336
rect 7872 1388 7924 1394
rect 7872 1330 7924 1336
rect 7976 1388 8028 1394
rect 7976 1330 8028 1336
rect 9645 1388 9697 1394
rect 9645 1330 9697 1336
rect 11290 1388 11342 1394
rect 11290 1330 11342 1336
rect 11472 1388 11524 1394
rect 11472 1330 11524 1336
rect 13036 1388 13088 1394
rect 13036 1330 13088 1336
rect 13223 1388 13275 1394
rect 13223 1330 13275 1336
rect 14880 1388 14932 1394
rect 14880 1330 14932 1336
rect 15159 1388 15211 1394
rect 15159 1330 15211 1336
rect 4673 1310 4737 1316
rect 4673 1258 4679 1310
rect 4731 1258 4737 1310
rect 4673 1252 4737 1258
rect 6421 1310 6485 1316
rect 6421 1258 6427 1310
rect 6479 1258 6485 1310
rect 9917 1310 9981 1316
rect 6421 1252 6485 1258
rect 8148 1293 8230 1299
rect 4031 928 4083 934
rect 4680 912 4730 1252
rect 5779 928 5831 934
rect 4031 870 4083 876
rect 4679 906 4731 912
rect 3719 699 3725 767
rect 3793 699 3799 767
rect 2261 314 2355 320
rect 4032 317 4081 870
rect 6428 912 6478 1252
rect 8148 1223 8154 1293
rect 8224 1223 8230 1293
rect 9917 1258 9923 1310
rect 9975 1258 9981 1310
rect 9917 1252 9981 1258
rect 11644 1293 11726 1299
rect 8148 1217 8230 1223
rect 7527 928 7579 934
rect 5779 870 5831 876
rect 6427 906 6479 912
rect 4679 848 4731 854
rect 5780 317 5829 870
rect 7527 870 7579 876
rect 8160 876 8218 1217
rect 6427 848 6479 854
rect 7528 317 7577 870
rect 9275 928 9327 934
rect 9924 912 9974 1252
rect 11644 1223 11650 1293
rect 11720 1223 11726 1293
rect 11644 1217 11726 1223
rect 13392 1293 13474 1299
rect 13392 1223 13398 1293
rect 13468 1223 13474 1293
rect 13392 1217 13474 1223
rect 11023 928 11075 934
rect 9275 870 9327 876
rect 9923 906 9975 912
rect 8160 812 8218 818
rect 9276 317 9325 870
rect 11023 870 11075 876
rect 11656 876 11714 1217
rect 9923 848 9975 854
rect 11024 317 11073 870
rect 12771 928 12823 934
rect 12771 870 12823 876
rect 13404 876 13462 1217
rect 15140 1208 15146 1260
rect 15198 1208 15204 1260
rect 11656 812 11714 818
rect 12772 317 12821 870
rect 14519 928 14571 934
rect 14519 870 14571 876
rect 15147 874 15197 1208
rect 13404 812 13462 818
rect 14520 317 14569 870
rect 15146 868 15198 874
rect 15146 810 15198 816
rect 60 307 119 313
rect 60 -139 119 248
rect 60 -204 119 -198
rect 1112 279 1164 285
rect 1112 221 1164 227
rect 2261 232 2267 314
rect 2349 232 2355 314
rect 4020 265 4026 317
rect 4087 265 4093 317
rect 5768 265 5774 317
rect 5835 265 5841 317
rect 7516 265 7522 317
rect 7583 265 7589 317
rect 9264 265 9270 317
rect 9331 265 9337 317
rect 11012 265 11018 317
rect 11079 265 11085 317
rect 12760 265 12766 317
rect 12827 265 12833 317
rect 14508 265 14514 317
rect 14575 265 14581 317
rect 2261 226 2355 232
rect 1112 -169 1163 221
rect 1112 -175 1164 -169
rect 1112 -233 1164 -227
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 28801
transform 1 0 47 0 -1 36
box -38 -48 406 592
use sky130_ef_sc_hd__fill_12  sky130_ef_sc_hd__fill_12_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 47 0 -1 1124
box -38 -48 1142 592
use sky130_ef_sc_hd__fill_12  sky130_ef_sc_hd__fill_12_1
timestamp 1646787781
transform 1 0 1151 0 -1 1124
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 2255 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_1
timestamp 1646787781
transform -1 0 1979 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_2
timestamp 1646787781
transform -1 0 1703 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_3
timestamp 1646787781
transform -1 0 1427 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_4
timestamp 1646787781
transform -1 0 2531 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_5
timestamp 1646787781
transform -1 0 4279 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_6
timestamp 1646787781
transform -1 0 6027 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_7
timestamp 1646787781
transform -1 0 7775 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_8
timestamp 1646787781
transform -1 0 9523 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_9
timestamp 1646787781
transform -1 0 11271 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_10
timestamp 1646787781
transform -1 0 13019 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_11
timestamp 1646787781
transform -1 0 14767 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 47 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1646787781
transform 1 0 323 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1646787781
transform 1 0 599 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1646787781
transform 1 0 875 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1646787781
transform -1 0 1151 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1646787781
transform -1 0 875 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1646787781
transform -1 0 599 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1646787781
transform 1 0 3727 0 -1 2212
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 4003 0 -1 2212
box -38 -48 682 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 2255 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1646787781
transform 1 0 4003 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1646787781
transform 1 0 5751 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1646787781
transform 1 0 7499 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4
timestamp 1646787781
transform 1 0 9247 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_5
timestamp 1646787781
transform 1 0 10995 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_6
timestamp 1646787781
transform 1 0 12743 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 4739 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_1
timestamp 1646787781
transform -1 0 6487 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_2
timestamp 1646787781
transform -1 0 8235 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_3
timestamp 1646787781
transform -1 0 9983 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_4
timestamp 1646787781
transform -1 0 11731 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_5
timestamp 1646787781
transform -1 0 13479 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_6
timestamp 1646787781
transform -1 0 15227 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  sky130_fd_sc_hd__einvn_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 3543 0 -1 1124
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 3543 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1646787781
transform 1 0 4739 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1646787781
transform 1 0 5475 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1646787781
transform 1 0 6487 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1646787781
transform 1 0 7223 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1646787781
transform 1 0 8235 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1646787781
transform 1 0 8971 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1646787781
transform 1 0 9983 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_9
timestamp 1646787781
transform 1 0 10719 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_10
timestamp 1646787781
transform 1 0 11731 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1646787781
transform 1 0 12467 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1646787781
transform 1 0 13479 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1646787781
transform 1 0 14215 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1646787781
transform 1 0 47 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1646787781
transform 1 0 783 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1646787781
transform 1 0 1519 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1646787781
transform 1 0 2255 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_18
timestamp 1646787781
transform 1 0 2991 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_19
timestamp 1646787781
transform 1 0 3727 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_20
timestamp 1646787781
transform 1 0 4739 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_21
timestamp 1646787781
transform 1 0 5475 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_22
timestamp 1646787781
transform 1 0 6487 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_23
timestamp 1646787781
transform 1 0 7223 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_24
timestamp 1646787781
transform 1 0 8235 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_25
timestamp 1646787781
transform 1 0 8971 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_26
timestamp 1646787781
transform 1 0 9983 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_27
timestamp 1646787781
transform 1 0 10719 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_28
timestamp 1646787781
transform 1 0 11731 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_29
timestamp 1646787781
transform 1 0 12467 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_30
timestamp 1646787781
transform 1 0 13479 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_31
timestamp 1646787781
transform 1 0 14215 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_32
timestamp 1646787781
transform 1 0 14491 0 1 36
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 14859 0 1 1124
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 7683 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_1
timestamp 1646787781
transform 1 0 11179 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_2
timestamp 1646787781
transform 1 0 12927 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  sky130_fd_sc_hd__or3_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 3083 0 1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 4095 0 1 1124
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_1
timestamp 1646787781
transform 1 0 5843 0 1 1124
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_2
timestamp 1646787781
transform 1 0 9339 0 1 1124
box -38 -48 682 592
<< labels >>
flabel metal1 s 47 1554 76 1583 1 FreeSerif 320 0 0 0 cfg_in[0]
flabel metal1 s 47 1486 76 1515 1 FreeSerif 320 0 0 0 cfg_in[1]
flabel metal1 s 47 1418 76 1447 1 FreeSerif 320 0 0 0 cfg_in[2]
<< end >>
