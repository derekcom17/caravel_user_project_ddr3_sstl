magic
tech sky130A
magscale 1 2
timestamp 1647071613
<< checkpaint >>
rect 8957 8368 18461 8912
rect 1413 6736 18461 8368
rect -243 5648 18461 6736
rect -3923 -3944 19197 5648
rect -3923 -4488 5213 -3944
<< nwell >>
rect 9929 3882 9945 4127
rect 9929 2794 9945 3039
rect 4685 1706 4885 1951
rect 9929 1706 9945 1951
<< psubdiff >>
rect 9880 4404 9931 4438
rect 9965 4404 10011 4438
rect 7081 -14 7132 20
rect 7166 -14 7212 20
rect 11900 -14 11951 20
rect 11985 -14 12031 20
<< psubdiffcont >>
rect 9931 4404 9965 4438
rect 7132 -14 7166 20
rect 11951 -14 11985 20
<< locali >>
rect 9880 4404 9931 4438
rect 9965 4404 10011 4438
rect 9891 4371 9983 4404
rect 14322 2923 14356 2960
rect 3749 2311 3790 2336
rect 3910 2004 3957 2031
rect 14322 1835 14356 1872
rect 2481 872 2637 913
rect 4228 861 4340 895
rect 5976 861 6088 895
rect 7724 861 7836 895
rect 9472 861 9584 895
rect 11220 861 11332 895
rect 12968 861 13080 895
rect 14716 861 14828 895
rect 4309 699 4388 767
rect 4456 699 4527 767
rect 2206 308 2343 361
rect 200 188 388 294
rect 476 188 665 294
rect 752 188 943 294
rect 1134 233 1172 307
rect 2206 291 2273 308
rect 1376 250 1497 284
rect 1652 253 1774 287
rect 1928 257 2053 291
rect 3938 262 4032 311
rect 5686 262 5780 311
rect 7434 262 7528 311
rect 9182 262 9276 311
rect 10930 262 11024 311
rect 12678 262 12772 311
rect 14426 262 14520 311
rect 2273 231 2343 238
rect 3940 247 3987 262
rect 3940 203 3941 247
rect 3985 203 3987 247
rect 3940 202 3987 203
rect 5688 247 5735 262
rect 5688 203 5689 247
rect 5733 203 5735 247
rect 5688 202 5735 203
rect 7436 247 7483 262
rect 7436 203 7437 247
rect 7481 203 7483 247
rect 7436 202 7483 203
rect 9184 247 9231 262
rect 9184 203 9185 247
rect 9229 203 9231 247
rect 9184 202 9231 203
rect 10932 247 10979 262
rect 10932 203 10933 247
rect 10977 203 10979 247
rect 10932 202 10979 203
rect 12680 247 12727 262
rect 12680 203 12681 247
rect 12725 203 12727 247
rect 12680 202 12727 203
rect 14428 247 14475 262
rect 14428 203 14429 247
rect 14473 203 14475 247
rect 14428 202 14475 203
rect 7081 -14 7132 20
rect 7166 -14 7212 20
rect 11900 -14 11951 20
rect 11985 -14 12031 20
rect 532 -222 722 -116
rect 809 -222 998 -116
<< viali >>
rect 14317 4620 14357 4660
rect 14070 4571 14110 4611
rect 12980 4484 13014 4518
rect 5749 4210 5805 4244
rect 6900 4210 6934 4244
rect 7237 4210 7271 4244
rect 8372 4210 8406 4244
rect 8709 4210 8743 4244
rect 9844 4210 9878 4244
rect 10273 4210 10307 4244
rect 11408 4210 11442 4244
rect 11745 4210 11779 4244
rect 12880 4210 12914 4244
rect 13217 4210 13251 4244
rect 5508 4130 5556 4178
rect 6994 4137 7028 4171
rect 8464 4137 8498 4171
rect 10026 4137 10060 4171
rect 11491 4137 11525 4171
rect 12963 4137 12997 4171
rect 14317 4011 14351 4045
rect 6877 3517 6911 3551
rect 8349 3517 8383 3551
rect 9814 3517 9848 3551
rect 11376 3517 11410 3551
rect 12846 3517 12880 3551
rect 14318 3510 14366 3558
rect 5515 3413 5559 3457
rect 6623 3444 6657 3478
rect 6960 3444 6994 3478
rect 8095 3444 8129 3478
rect 8432 3444 8466 3478
rect 9567 3444 9601 3478
rect 11131 3444 11165 3478
rect 11468 3444 11502 3478
rect 12603 3444 12637 3478
rect 12940 3444 12974 3478
rect 14071 3445 14114 3479
rect 10029 3406 10063 3440
rect 5749 3122 5805 3156
rect 6900 3122 6934 3156
rect 7237 3122 7271 3156
rect 8372 3122 8406 3156
rect 8709 3122 8743 3156
rect 9844 3122 9878 3156
rect 10273 3122 10307 3156
rect 11408 3122 11442 3156
rect 11745 3122 11779 3156
rect 12880 3122 12914 3156
rect 13217 3122 13251 3156
rect 5508 3042 5556 3090
rect 6994 3049 7028 3083
rect 8464 3049 8498 3083
rect 10026 3049 10060 3083
rect 11491 3049 11525 3083
rect 12963 3049 12997 3083
rect 14322 2960 14356 2994
rect 5135 2501 5169 2535
rect 4138 2427 4172 2461
rect 5256 2438 5296 2472
rect 6877 2429 6911 2463
rect 8349 2429 8383 2463
rect 9814 2429 9848 2463
rect 11376 2429 11410 2463
rect 12846 2429 12880 2463
rect 14318 2422 14366 2470
rect 3749 2336 3790 2377
rect 5515 2325 5559 2369
rect 6623 2356 6657 2390
rect 6960 2356 6994 2390
rect 8095 2356 8129 2390
rect 8432 2356 8466 2390
rect 9567 2356 9601 2390
rect 10029 2325 10063 2359
rect 11131 2356 11165 2390
rect 11468 2356 11502 2390
rect 12603 2356 12637 2390
rect 12940 2356 12974 2390
rect 14071 2357 14114 2391
rect 6820 2034 6854 2068
rect 7236 2034 7270 2068
rect 8372 2034 8406 2068
rect 8709 2034 8743 2068
rect 9844 2034 9878 2068
rect 10273 2034 10307 2068
rect 11408 2034 11442 2068
rect 11745 2034 11779 2068
rect 12880 2034 12914 2068
rect 13217 2034 13251 2068
rect 3731 1978 3787 2034
rect 3910 1957 3957 2004
rect 4119 1963 4154 1998
rect 4570 1948 4630 2008
rect 5044 1954 5092 2002
rect 5387 1954 5427 1994
rect 6994 1961 7028 1995
rect 8464 1961 8498 1995
rect 10026 1961 10060 1995
rect 11491 1961 11525 1995
rect 12963 1961 12997 1995
rect 14322 1872 14356 1906
rect 6821 1753 6855 1787
rect 3288 1549 3322 1583
rect 4313 1549 4347 1583
rect 6057 1549 6091 1583
rect 9468 1549 9502 1583
rect 3207 1413 3241 1447
rect 4400 1413 4434 1447
rect 6148 1413 6182 1447
rect 3115 1324 3155 1364
rect 4120 1342 4160 1382
rect 5878 1342 5918 1382
rect 7792 1345 7826 1379
rect 7878 1342 7918 1382
rect 7982 1342 8022 1382
rect 9370 1345 9404 1379
rect 9651 1342 9691 1382
rect 11296 1342 11336 1382
rect 11384 1345 11418 1379
rect 11478 1342 11518 1382
rect 13042 1342 13082 1382
rect 13138 1345 13172 1379
rect 13229 1342 13269 1382
rect 14886 1342 14926 1382
rect 15038 1345 15072 1379
rect 15165 1342 15205 1382
rect 3491 1261 3525 1295
rect 4688 1267 4722 1301
rect 6436 1267 6470 1301
rect 8160 1229 8218 1287
rect 9932 1267 9966 1301
rect 11656 1229 11714 1287
rect 13404 1229 13462 1287
rect 15155 1217 15189 1251
rect 2279 867 2337 925
rect 2749 888 2805 944
rect 3488 876 3528 916
rect 4037 882 4077 922
rect 4685 860 4725 900
rect 5785 882 5825 922
rect 6433 860 6473 900
rect 7533 882 7573 922
rect 9281 882 9321 922
rect 8166 824 8212 870
rect 9929 860 9969 900
rect 11029 882 11069 922
rect 12777 882 12817 922
rect 11662 824 11708 870
rect 14525 882 14565 922
rect 13410 824 13456 870
rect 15152 822 15192 862
rect 4388 699 4456 767
rect 6135 705 6191 761
rect 7922 705 7978 761
rect 9641 705 9697 761
rect 11372 705 11428 761
rect 13127 705 13183 761
rect 14884 705 14940 761
rect 66 254 113 301
rect 1060 234 1099 273
rect 2273 238 2343 308
rect 4032 262 4081 311
rect 5780 262 5829 311
rect 7528 262 7577 311
rect 9276 262 9325 311
rect 11024 262 11073 311
rect 12772 262 12821 311
rect 14520 262 14569 311
rect 2529 197 2585 253
rect 3941 203 3985 247
rect 4277 197 4333 253
rect 5689 203 5733 247
rect 6025 197 6081 253
rect 7437 203 7481 247
rect 7773 197 7829 253
rect 9185 203 9229 247
rect 9521 197 9577 253
rect 10933 203 10977 247
rect 11269 197 11325 253
rect 12681 203 12725 247
rect 13017 197 13073 253
rect 14429 203 14473 247
rect 344 -222 403 -116
rect 1118 -221 1158 -181
<< metal1 >>
rect 4123 4566 4129 4618
rect 4181 4602 4187 4618
rect 11387 4602 11393 4614
rect 4181 4574 11393 4602
rect 4181 4566 4187 4574
rect 11387 4562 11393 4574
rect 11445 4562 11451 4614
rect 14058 4565 14064 4617
rect 14116 4565 14122 4617
rect 14305 4614 14311 4666
rect 14363 4614 14369 4666
rect 5120 4472 5126 4524
rect 5178 4518 5184 4524
rect 12974 4518 13026 4524
rect 5178 4484 12980 4518
rect 13014 4484 13026 4518
rect 5178 4472 5184 4484
rect 12974 4478 13026 4484
rect 9891 4340 9983 4436
rect 11393 4279 11445 4285
rect 5743 4250 5749 4260
rect 5737 4204 5749 4250
rect 5805 4250 5811 4260
rect 5805 4204 5817 4250
rect 6888 4244 6946 4250
rect 6888 4210 6900 4244
rect 6934 4241 6946 4244
rect 7225 4244 7283 4250
rect 7225 4241 7237 4244
rect 6934 4213 7237 4241
rect 6934 4210 6946 4213
rect 6888 4204 6946 4210
rect 7225 4210 7237 4213
rect 7271 4210 7283 4244
rect 7225 4204 7283 4210
rect 8360 4244 8418 4250
rect 8360 4210 8372 4244
rect 8406 4241 8418 4244
rect 8697 4244 8755 4250
rect 8697 4241 8709 4244
rect 8406 4213 8709 4241
rect 8406 4210 8418 4213
rect 8360 4204 8418 4210
rect 8697 4210 8709 4213
rect 8743 4210 8755 4244
rect 8697 4204 8755 4210
rect 9832 4244 9890 4250
rect 9832 4210 9844 4244
rect 9878 4241 9890 4244
rect 10261 4244 10319 4250
rect 10261 4241 10273 4244
rect 9878 4213 10273 4241
rect 9878 4210 9890 4213
rect 9832 4204 9890 4210
rect 10261 4210 10273 4213
rect 10307 4210 10319 4244
rect 11445 4241 11454 4250
rect 11733 4244 11791 4250
rect 11733 4241 11745 4244
rect 11445 4227 11745 4241
rect 11393 4221 11408 4227
rect 10261 4204 10319 4210
rect 11396 4210 11408 4221
rect 11442 4213 11745 4227
rect 11442 4210 11454 4213
rect 11396 4204 11454 4210
rect 11733 4210 11745 4213
rect 11779 4210 11791 4244
rect 11733 4204 11791 4210
rect 12868 4244 12926 4250
rect 12868 4210 12880 4244
rect 12914 4241 12926 4244
rect 13205 4244 13263 4250
rect 13205 4241 13217 4244
rect 12914 4213 13217 4241
rect 12914 4210 12926 4213
rect 12868 4204 12926 4210
rect 13205 4210 13217 4213
rect 13251 4210 13263 4244
rect 13205 4204 13263 4210
rect 5495 4184 5501 4188
rect 5437 4136 5501 4184
rect 5553 4184 5559 4188
rect 5553 4178 5568 4184
rect 5556 4175 5568 4178
rect 6982 4175 7040 4177
rect 8458 4175 8504 4183
rect 10014 4175 10072 4177
rect 11479 4175 11537 4177
rect 12957 4175 13003 4183
rect 14305 4175 14311 4180
rect 5556 4171 14311 4175
rect 5556 4137 6994 4171
rect 7028 4137 8464 4171
rect 8498 4137 10026 4171
rect 10060 4137 11491 4171
rect 11525 4137 12963 4171
rect 12997 4137 14311 4171
rect 5437 4130 5508 4136
rect 5556 4133 14311 4137
rect 5556 4130 5568 4133
rect 6982 4131 7040 4133
rect 5437 4124 5568 4130
rect 8458 4125 8504 4133
rect 10014 4131 10072 4133
rect 11479 4131 11537 4133
rect 12957 4125 13003 4133
rect 14305 4128 14311 4133
rect 14363 4128 14369 4180
rect 14058 4002 14064 4054
rect 14116 4045 14122 4054
rect 14305 4045 14363 4051
rect 14116 4011 14317 4045
rect 14351 4011 14363 4045
rect 14116 4002 14122 4011
rect 14305 4005 14363 4011
rect 5495 3508 5501 3560
rect 5553 3555 5559 3560
rect 6871 3555 6917 3563
rect 8337 3555 8395 3557
rect 9802 3555 9860 3557
rect 11370 3555 11416 3563
rect 12834 3555 12892 3557
rect 14302 3555 14308 3567
rect 14360 3564 14366 3567
rect 14360 3558 14437 3564
rect 5553 3551 14308 3555
rect 5553 3517 6877 3551
rect 6911 3517 8349 3551
rect 8383 3517 9814 3551
rect 9848 3517 11376 3551
rect 11410 3517 12846 3551
rect 12880 3517 14308 3551
rect 5553 3515 14308 3517
rect 5553 3513 14318 3515
rect 5553 3508 5559 3513
rect 6871 3505 6917 3513
rect 8337 3511 8395 3513
rect 9802 3511 9860 3513
rect 11370 3505 11416 3513
rect 12834 3511 12892 3513
rect 14306 3510 14318 3513
rect 14366 3510 14437 3558
rect 14306 3504 14437 3510
rect 6611 3478 6669 3484
rect 5503 3457 5749 3463
rect 5503 3413 5515 3457
rect 5559 3413 5749 3457
rect 5503 3407 5749 3413
rect 5805 3407 5811 3463
rect 6611 3444 6623 3478
rect 6657 3475 6669 3478
rect 6948 3478 7006 3484
rect 6948 3475 6960 3478
rect 6657 3447 6960 3475
rect 6657 3444 6669 3447
rect 6611 3438 6669 3444
rect 6948 3444 6960 3447
rect 6994 3444 7006 3478
rect 6948 3438 7006 3444
rect 8083 3478 8141 3484
rect 8083 3444 8095 3478
rect 8129 3475 8141 3478
rect 8420 3478 8478 3484
rect 8420 3475 8432 3478
rect 8129 3447 8432 3475
rect 8129 3444 8141 3447
rect 8083 3438 8141 3444
rect 8420 3444 8432 3447
rect 8466 3444 8478 3478
rect 8420 3438 8478 3444
rect 9555 3478 9613 3484
rect 9555 3444 9567 3478
rect 9601 3475 9613 3478
rect 11119 3478 11177 3484
rect 9601 3452 10060 3475
rect 9601 3447 10069 3452
rect 9601 3444 9613 3447
rect 9555 3438 9613 3444
rect 10023 3440 10069 3447
rect 10023 3406 10029 3440
rect 10063 3406 10069 3440
rect 11119 3444 11131 3478
rect 11165 3475 11177 3478
rect 11456 3478 11514 3484
rect 11456 3475 11468 3478
rect 11165 3447 11468 3475
rect 11165 3444 11177 3447
rect 11119 3438 11177 3444
rect 11456 3444 11468 3447
rect 11502 3444 11514 3478
rect 11456 3438 11514 3444
rect 12591 3478 12649 3484
rect 12591 3444 12603 3478
rect 12637 3475 12649 3478
rect 12928 3478 12986 3484
rect 12928 3475 12940 3478
rect 12637 3447 12940 3475
rect 12637 3444 12649 3447
rect 12591 3438 12649 3444
rect 12928 3444 12940 3447
rect 12974 3444 12986 3478
rect 12928 3438 12986 3444
rect 14059 3433 14068 3485
rect 14120 3433 14126 3485
rect 10023 3394 10069 3406
rect 5743 3162 5749 3172
rect 5737 3116 5749 3162
rect 5805 3162 5811 3172
rect 5805 3116 5817 3162
rect 6888 3156 6946 3162
rect 6888 3122 6900 3156
rect 6934 3153 6946 3156
rect 7225 3156 7283 3162
rect 7225 3153 7237 3156
rect 6934 3125 7237 3153
rect 6934 3122 6946 3125
rect 6888 3116 6946 3122
rect 7225 3122 7237 3125
rect 7271 3122 7283 3156
rect 7225 3116 7283 3122
rect 8360 3156 8418 3162
rect 8360 3122 8372 3156
rect 8406 3153 8418 3156
rect 8697 3156 8755 3162
rect 8697 3153 8709 3156
rect 8406 3125 8709 3153
rect 8406 3122 8418 3125
rect 8360 3116 8418 3122
rect 8697 3122 8709 3125
rect 8743 3122 8755 3156
rect 8697 3116 8755 3122
rect 9832 3156 9890 3162
rect 9832 3122 9844 3156
rect 9878 3153 9890 3156
rect 10261 3156 10319 3162
rect 10261 3153 10273 3156
rect 9878 3125 10273 3153
rect 9878 3122 9890 3125
rect 9832 3116 9890 3122
rect 10261 3122 10273 3125
rect 10307 3122 10319 3156
rect 10261 3116 10319 3122
rect 11396 3156 11454 3162
rect 11396 3122 11408 3156
rect 11442 3153 11454 3156
rect 11733 3156 11791 3162
rect 11733 3153 11745 3156
rect 11442 3125 11745 3153
rect 11442 3122 11454 3125
rect 11396 3116 11454 3122
rect 11733 3122 11745 3125
rect 11779 3122 11791 3156
rect 11733 3116 11791 3122
rect 12868 3156 12926 3162
rect 12868 3122 12880 3156
rect 12914 3153 12926 3156
rect 13205 3156 13263 3162
rect 13205 3153 13217 3156
rect 12914 3125 13217 3153
rect 12914 3122 12926 3125
rect 12868 3116 12926 3122
rect 13205 3122 13217 3125
rect 13251 3122 13263 3156
rect 13205 3116 13263 3122
rect 5504 3096 5510 3100
rect 5437 3090 5510 3096
rect 5437 3042 5508 3090
rect 5562 3087 5568 3100
rect 6982 3087 7040 3089
rect 8458 3087 8504 3095
rect 10014 3087 10072 3089
rect 11479 3087 11537 3089
rect 12957 3087 13003 3095
rect 14302 3087 14308 3092
rect 5562 3083 14308 3087
rect 5562 3049 6994 3083
rect 7028 3049 8464 3083
rect 8498 3049 10026 3083
rect 10060 3049 11491 3083
rect 11525 3049 12963 3083
rect 12997 3049 14308 3083
rect 5562 3048 14308 3049
rect 5556 3045 14308 3048
rect 5556 3042 5568 3045
rect 6982 3043 7040 3045
rect 5437 3036 5568 3042
rect 8458 3037 8504 3045
rect 10014 3043 10072 3045
rect 11479 3043 11537 3045
rect 12957 3037 13003 3045
rect 14302 3040 14308 3045
rect 14360 3040 14366 3092
rect 14062 2951 14068 3003
rect 14120 2994 14126 3003
rect 14310 2994 14368 3000
rect 14120 2960 14322 2994
rect 14356 2960 14368 2994
rect 14120 2951 14126 2960
rect 14310 2954 14368 2960
rect 5881 2665 5887 2677
rect 3587 2637 5887 2665
rect 5881 2625 5887 2637
rect 5939 2625 5945 2677
rect 5120 2492 5126 2544
rect 5178 2492 5184 2544
rect 4123 2470 4187 2476
rect 4123 2418 4129 2470
rect 4181 2418 4187 2470
rect 5244 2432 5250 2484
rect 5302 2432 5308 2484
rect 14316 2476 14322 2478
rect 5250 2426 5302 2432
rect 5504 2420 5510 2472
rect 5562 2467 5568 2472
rect 6871 2467 6917 2475
rect 8337 2467 8395 2469
rect 9802 2467 9860 2469
rect 11370 2467 11416 2475
rect 14306 2470 14322 2476
rect 14374 2476 14380 2478
rect 12834 2467 12892 2469
rect 14306 2467 14318 2470
rect 5562 2463 14318 2467
rect 5562 2429 6877 2463
rect 6911 2429 8349 2463
rect 8383 2429 9814 2463
rect 9848 2429 11376 2463
rect 11410 2429 12846 2463
rect 12880 2429 14318 2463
rect 5562 2425 14318 2429
rect 14374 2426 14437 2476
rect 5562 2420 5568 2425
rect 4123 2412 4187 2418
rect 6871 2417 6917 2425
rect 8337 2423 8395 2425
rect 9802 2423 9860 2425
rect 11370 2417 11416 2425
rect 12834 2423 12892 2425
rect 14306 2422 14318 2425
rect 14366 2422 14437 2426
rect 14306 2416 14437 2422
rect 6611 2390 6669 2396
rect 3737 2377 3802 2383
rect 4464 2377 4470 2383
rect 3586 2336 3749 2377
rect 3790 2336 4470 2377
rect 3737 2330 3802 2336
rect 4464 2331 4470 2336
rect 4522 2331 4528 2383
rect 5503 2369 5749 2375
rect 5503 2325 5515 2369
rect 5559 2325 5749 2369
rect 5503 2319 5749 2325
rect 5805 2319 5811 2375
rect 6611 2356 6623 2390
rect 6657 2387 6669 2390
rect 6948 2390 7006 2396
rect 6948 2387 6960 2390
rect 6657 2359 6960 2387
rect 6657 2356 6669 2359
rect 6611 2350 6669 2356
rect 6948 2356 6960 2359
rect 6994 2356 7006 2390
rect 6948 2350 7006 2356
rect 8083 2390 8141 2396
rect 8083 2356 8095 2390
rect 8129 2387 8141 2390
rect 8420 2390 8478 2396
rect 8420 2387 8432 2390
rect 8129 2359 8432 2387
rect 8129 2356 8141 2359
rect 8083 2350 8141 2356
rect 8420 2356 8432 2359
rect 8466 2356 8478 2390
rect 8420 2350 8478 2356
rect 9555 2390 9613 2396
rect 9555 2356 9567 2390
rect 9601 2387 9613 2390
rect 11119 2390 11177 2396
rect 9601 2371 10060 2387
rect 9601 2359 10069 2371
rect 9601 2356 9613 2359
rect 9555 2350 9613 2356
rect 10023 2325 10029 2359
rect 10063 2325 10069 2359
rect 11119 2356 11131 2390
rect 11165 2387 11177 2390
rect 11456 2390 11514 2396
rect 11456 2387 11468 2390
rect 11165 2359 11468 2387
rect 11165 2356 11177 2359
rect 11119 2350 11177 2356
rect 11456 2356 11468 2359
rect 11502 2356 11514 2390
rect 11456 2350 11514 2356
rect 12591 2390 12649 2396
rect 12591 2356 12603 2390
rect 12637 2387 12649 2390
rect 12928 2390 12986 2396
rect 12928 2387 12940 2390
rect 12637 2359 12940 2387
rect 12637 2356 12649 2359
rect 12591 2350 12649 2356
rect 12928 2356 12940 2359
rect 12974 2356 12986 2390
rect 12928 2350 12986 2356
rect 14059 2345 14068 2397
rect 14120 2345 14126 2397
rect 10023 2313 10069 2325
rect 4465 2082 4471 2134
rect 4523 2129 4529 2134
rect 4523 2124 5193 2129
rect 5375 2124 5381 2136
rect 4523 2096 5381 2124
rect 4523 2088 5193 2096
rect 4523 2082 4529 2088
rect 5375 2084 5381 2096
rect 5433 2084 5439 2136
rect 6808 2068 6866 2074
rect 3719 1972 3725 2040
rect 3793 1972 3799 2040
rect 3898 2004 3969 2010
rect 4564 2008 4636 2020
rect 5881 2016 5887 2068
rect 5939 2016 5945 2068
rect 6808 2034 6820 2068
rect 6854 2065 6866 2068
rect 7224 2068 7283 2074
rect 7224 2065 7236 2068
rect 6854 2037 7236 2065
rect 6854 2034 6866 2037
rect 6808 2028 6866 2034
rect 7224 2034 7236 2037
rect 7270 2034 7283 2068
rect 7224 2028 7283 2034
rect 8360 2068 8418 2074
rect 8360 2034 8372 2068
rect 8406 2065 8418 2068
rect 8697 2068 8755 2074
rect 8697 2065 8709 2068
rect 8406 2037 8709 2065
rect 8406 2034 8418 2037
rect 8360 2028 8418 2034
rect 8697 2034 8709 2037
rect 8743 2034 8755 2068
rect 8697 2028 8755 2034
rect 9832 2068 9890 2074
rect 9832 2034 9844 2068
rect 9878 2065 9890 2068
rect 10261 2068 10319 2074
rect 10261 2065 10273 2068
rect 9878 2037 10273 2065
rect 9878 2034 9890 2037
rect 9832 2028 9890 2034
rect 10261 2034 10273 2037
rect 10307 2034 10319 2068
rect 10261 2028 10319 2034
rect 11396 2068 11454 2074
rect 11396 2034 11408 2068
rect 11442 2065 11454 2068
rect 11733 2068 11791 2074
rect 11733 2065 11745 2068
rect 11442 2037 11745 2065
rect 11442 2034 11454 2037
rect 11396 2028 11454 2034
rect 11733 2034 11745 2037
rect 11779 2034 11791 2068
rect 11733 2028 11791 2034
rect 12868 2068 12926 2074
rect 12868 2034 12880 2068
rect 12914 2065 12926 2068
rect 13205 2068 13263 2074
rect 13205 2065 13217 2068
rect 12914 2037 13217 2065
rect 12914 2034 12926 2037
rect 12868 2028 12926 2034
rect 13205 2034 13217 2037
rect 13251 2034 13263 2068
rect 13205 2028 13263 2034
rect 3898 1957 3910 2004
rect 3957 1998 4166 2004
rect 3957 1963 4119 1998
rect 4154 1963 4166 1998
rect 3957 1957 4166 1963
rect 3898 1951 3969 1957
rect 4564 1948 4570 2008
rect 4630 2002 5104 2008
rect 4630 1954 5044 2002
rect 5092 1986 5104 2002
rect 5092 1958 5166 1986
rect 5092 1954 5104 1958
rect 4630 1948 5104 1954
rect 4564 1936 4636 1948
rect 5138 1920 5166 1958
rect 5375 1948 5381 2000
rect 5433 1948 5439 2000
rect 6982 1999 7040 2001
rect 8458 1999 8504 2007
rect 10014 1999 10072 2001
rect 11479 1999 11537 2001
rect 12957 1999 13003 2007
rect 14316 1999 14322 2004
rect 6976 1995 14322 1999
rect 6976 1990 6994 1995
rect 6890 1962 6994 1990
rect 6890 1920 6918 1962
rect 6976 1961 6994 1962
rect 7028 1961 8464 1995
rect 8498 1961 10026 1995
rect 10060 1961 11491 1995
rect 11525 1961 12963 1995
rect 12997 1961 14322 1995
rect 6976 1957 14322 1961
rect 6982 1955 7040 1957
rect 8458 1949 8504 1957
rect 10014 1955 10072 1957
rect 11479 1955 11537 1957
rect 12957 1949 13003 1957
rect 14316 1952 14322 1957
rect 14374 1952 14380 2004
rect 5138 1892 6918 1920
rect 14062 1863 14068 1915
rect 14120 1906 14126 1915
rect 14310 1906 14368 1912
rect 14120 1872 14322 1906
rect 14356 1872 14368 1906
rect 14120 1863 14126 1872
rect 14310 1866 14368 1872
rect 5238 1784 5244 1796
rect 5226 1756 5244 1784
rect 5238 1744 5244 1756
rect 5296 1784 5302 1796
rect 6809 1787 6867 1793
rect 6809 1784 6821 1787
rect 5296 1756 6821 1784
rect 5296 1744 5302 1756
rect 6809 1753 6821 1756
rect 6855 1753 6867 1787
rect 6809 1747 6867 1753
rect 3276 1583 3334 1589
rect 4108 1583 4114 1592
rect 47 1552 3288 1583
rect 47 1549 3081 1552
rect 3189 1549 3288 1552
rect 3322 1549 4114 1583
rect 3276 1543 3334 1549
rect 4108 1540 4114 1549
rect 4166 1540 4172 1592
rect 4301 1583 4359 1592
rect 4301 1549 4313 1583
rect 4347 1549 4359 1583
rect 3103 1515 3109 1524
rect 47 1481 3109 1515
rect 3103 1472 3109 1481
rect 3161 1515 3167 1524
rect 4301 1515 4359 1549
rect 4485 1540 4491 1592
rect 4543 1583 4549 1592
rect 6045 1583 6103 1589
rect 7970 1583 7976 1592
rect 4543 1552 6057 1583
rect 4543 1549 5838 1552
rect 5958 1549 6057 1552
rect 6091 1552 7976 1583
rect 6091 1549 7844 1552
rect 7952 1549 7976 1552
rect 4543 1540 4549 1549
rect 6045 1543 6103 1549
rect 7970 1540 7976 1549
rect 8028 1583 8034 1592
rect 9462 1583 9508 1589
rect 11466 1583 11472 1592
rect 8028 1549 9468 1583
rect 9502 1552 11472 1583
rect 9502 1549 9617 1552
rect 9725 1549 11256 1552
rect 11376 1549 11472 1552
rect 8028 1540 8034 1549
rect 9462 1543 9508 1549
rect 11466 1540 11472 1549
rect 11524 1583 11530 1592
rect 13030 1583 13036 1592
rect 11524 1549 13036 1583
rect 11524 1540 11530 1549
rect 13030 1540 13036 1549
rect 13088 1583 13094 1592
rect 15153 1583 15159 1592
rect 13088 1552 15159 1583
rect 13088 1549 13195 1552
rect 13303 1549 14852 1552
rect 14960 1549 15159 1552
rect 13088 1540 13094 1549
rect 15153 1540 15159 1549
rect 15211 1583 15217 1592
rect 15211 1549 15227 1583
rect 15211 1540 15217 1549
rect 5866 1515 5872 1524
rect 3161 1512 4080 1515
rect 4200 1512 4457 1515
rect 4577 1512 5872 1515
rect 3161 1481 5872 1512
rect 3161 1472 3167 1481
rect 5866 1472 5872 1481
rect 5924 1515 5930 1524
rect 7866 1515 7872 1524
rect 5924 1481 7872 1515
rect 5924 1472 5930 1481
rect 7866 1472 7872 1481
rect 7924 1515 7930 1524
rect 9639 1515 9645 1524
rect 7924 1512 7942 1515
rect 8062 1512 9645 1515
rect 7924 1481 9645 1512
rect 7924 1472 7930 1481
rect 9639 1472 9645 1481
rect 9697 1515 9703 1524
rect 11284 1515 11290 1524
rect 9697 1481 11290 1515
rect 9697 1472 9703 1481
rect 11284 1472 11290 1481
rect 11342 1515 11348 1524
rect 13217 1515 13223 1524
rect 11342 1512 11444 1515
rect 11564 1512 13008 1515
rect 13116 1512 13223 1515
rect 11342 1481 13223 1512
rect 11342 1472 11348 1481
rect 13217 1472 13223 1481
rect 13275 1515 13281 1524
rect 14874 1515 14880 1524
rect 13275 1481 14880 1515
rect 13275 1472 13281 1481
rect 14874 1472 14880 1481
rect 14932 1515 14938 1524
rect 14932 1512 15131 1515
rect 14932 1481 15227 1512
rect 14932 1472 14938 1481
rect 3195 1447 3253 1453
rect 4388 1447 4446 1453
rect 6136 1447 6194 1453
rect 47 1444 3081 1447
rect 3189 1444 3207 1447
rect 47 1413 3207 1444
rect 3241 1416 4400 1447
rect 3241 1413 4080 1416
rect 4200 1413 4400 1416
rect 4434 1444 5838 1447
rect 5958 1444 6148 1447
rect 4434 1416 6148 1444
rect 4434 1413 5838 1416
rect 5958 1413 6148 1416
rect 6182 1444 7844 1447
rect 7964 1444 9617 1447
rect 9725 1444 11256 1447
rect 11376 1444 13195 1447
rect 13303 1444 14852 1447
rect 14960 1444 15227 1447
rect 6182 1416 15227 1444
rect 6182 1413 7838 1416
rect 8062 1413 9611 1416
rect 9731 1413 11256 1416
rect 11376 1413 11438 1416
rect 11558 1413 13002 1416
rect 13110 1413 13201 1416
rect 13309 1413 14846 1416
rect 14966 1413 15125 1416
rect 3195 1407 3253 1413
rect 4388 1407 4446 1413
rect 6136 1407 6194 1413
rect 3103 1318 3109 1370
rect 3161 1318 3167 1370
rect 4108 1333 4114 1388
rect 4166 1376 4172 1388
rect 4485 1376 4491 1385
rect 4166 1342 4491 1376
rect 4166 1333 4172 1342
rect 4485 1333 4491 1342
rect 4543 1333 4549 1385
rect 5866 1336 5872 1388
rect 5924 1336 5930 1388
rect 7786 1379 7832 1413
rect 7786 1345 7792 1379
rect 7826 1345 7832 1379
rect 7786 1333 7832 1345
rect 7866 1336 7872 1388
rect 7924 1336 7930 1388
rect 7970 1336 7976 1388
rect 8028 1336 8034 1388
rect 9364 1379 9410 1413
rect 9364 1345 9370 1379
rect 9404 1345 9410 1379
rect 9364 1333 9410 1345
rect 9639 1336 9645 1388
rect 9697 1336 9703 1388
rect 11284 1336 11290 1388
rect 11342 1336 11348 1388
rect 11378 1379 11424 1413
rect 11378 1345 11384 1379
rect 11418 1345 11424 1379
rect 11378 1333 11424 1345
rect 11466 1336 11472 1388
rect 11524 1336 11530 1388
rect 13030 1336 13036 1388
rect 13088 1336 13094 1388
rect 13132 1379 13178 1413
rect 13132 1345 13138 1379
rect 13172 1345 13178 1379
rect 13132 1333 13178 1345
rect 13217 1336 13223 1388
rect 13275 1336 13281 1388
rect 14874 1336 14880 1388
rect 14932 1336 14938 1388
rect 15032 1379 15078 1413
rect 15032 1345 15038 1379
rect 15072 1345 15078 1379
rect 15032 1333 15078 1345
rect 15153 1336 15159 1388
rect 15211 1336 15217 1388
rect 4679 1310 4731 1316
rect 3482 1304 3534 1310
rect 4679 1252 4731 1258
rect 6427 1310 6479 1316
rect 9923 1310 9975 1316
rect 6427 1252 6479 1258
rect 8148 1293 8230 1299
rect 3482 1246 3534 1252
rect 8148 1223 8154 1293
rect 8224 1223 8230 1293
rect 9923 1252 9975 1258
rect 11644 1293 11726 1299
rect 8148 1217 8230 1223
rect 11644 1223 11650 1293
rect 11720 1223 11726 1293
rect 11644 1217 11726 1223
rect 13392 1293 13474 1299
rect 13392 1223 13398 1293
rect 13468 1223 13474 1293
rect 13392 1217 13474 1223
rect 15146 1260 15198 1266
rect 15146 1202 15198 1208
rect 2743 944 2811 956
rect 2267 861 2273 931
rect 2343 861 2349 931
rect 2743 888 2749 944
rect 2805 888 2811 944
rect 2743 767 2811 888
rect 3476 870 3482 922
rect 3534 870 3540 922
rect 4025 876 4031 928
rect 4083 876 4089 928
rect 4673 854 4679 906
rect 4731 854 4737 906
rect 5773 876 5779 928
rect 5831 876 5837 928
rect 6421 854 6427 906
rect 6479 854 6485 906
rect 7521 876 7527 928
rect 7579 876 7585 928
rect 9269 876 9275 928
rect 9327 876 9333 928
rect 8154 818 8160 876
rect 8218 818 8224 876
rect 9917 854 9923 906
rect 9975 854 9981 906
rect 11017 876 11023 928
rect 11075 876 11081 928
rect 12765 876 12771 928
rect 12823 876 12829 928
rect 14513 876 14519 928
rect 14571 876 14577 928
rect 11650 818 11656 876
rect 11714 818 11720 876
rect 13398 818 13404 876
rect 13462 818 13468 876
rect 15140 816 15146 868
rect 15198 816 15204 868
rect 3725 767 3793 773
rect 4382 767 4462 779
rect 2743 699 3725 767
rect 3793 699 4388 767
rect 4456 761 15019 767
rect 4456 705 6135 761
rect 6191 705 7922 761
rect 7978 705 9641 761
rect 9697 705 11372 761
rect 11428 705 13127 761
rect 13183 705 14884 761
rect 14940 705 15019 761
rect 4456 699 15019 705
rect 3725 693 3793 699
rect 4382 687 4462 699
rect 2261 314 2355 320
rect 54 248 60 307
rect 119 248 125 307
rect 1048 273 1112 279
rect 1048 234 1060 273
rect 1099 234 1112 273
rect 1048 228 1112 234
rect 1106 227 1112 228
rect 1164 227 1170 279
rect 2261 232 2267 314
rect 2349 232 2355 314
rect 4026 317 4087 323
rect 5774 317 5835 323
rect 7522 317 7583 323
rect 9270 317 9331 323
rect 11018 317 11079 323
rect 12766 317 12827 323
rect 14514 317 14575 323
rect 2261 226 2355 232
rect 2523 253 2591 265
rect 4026 262 4032 265
rect 4081 262 4087 265
rect 2523 197 2529 253
rect 2585 247 3997 253
rect 4026 250 4087 262
rect 4271 253 4339 265
rect 5774 262 5780 265
rect 5829 262 5835 265
rect 2585 203 3941 247
rect 3985 203 3997 247
rect 2585 197 3997 203
rect 4271 197 4277 253
rect 4333 247 5745 253
rect 5774 250 5835 262
rect 6019 253 6087 265
rect 7522 262 7528 265
rect 7577 262 7583 265
rect 4333 203 5689 247
rect 5733 203 5745 247
rect 4333 197 5745 203
rect 6019 197 6025 253
rect 6081 247 7493 253
rect 7522 250 7583 262
rect 7767 253 7835 265
rect 9270 262 9276 265
rect 9325 262 9331 265
rect 6081 203 7437 247
rect 7481 203 7493 247
rect 6081 197 7493 203
rect 7767 197 7773 253
rect 7829 247 9241 253
rect 9270 250 9331 262
rect 9515 253 9583 265
rect 11018 262 11024 265
rect 11073 262 11079 265
rect 7829 203 9185 247
rect 9229 203 9241 247
rect 7829 197 9241 203
rect 9515 197 9521 253
rect 9577 247 10989 253
rect 11018 250 11079 262
rect 11263 253 11331 265
rect 12766 262 12772 265
rect 12821 262 12827 265
rect 9577 203 10933 247
rect 10977 203 10989 247
rect 9577 197 10989 203
rect 11263 197 11269 253
rect 11325 247 12737 253
rect 12766 250 12827 262
rect 13011 253 13079 265
rect 14514 262 14520 265
rect 14569 262 14575 265
rect 11325 203 12681 247
rect 12725 203 12737 247
rect 11325 197 12737 203
rect 13011 197 13017 253
rect 13073 247 14485 253
rect 14514 250 14575 262
rect 13073 203 14429 247
rect 14473 203 14485 247
rect 13073 197 14485 203
rect 2523 185 2591 197
rect 4271 185 4339 197
rect 6019 185 6087 197
rect 7767 185 7835 197
rect 9515 185 9583 197
rect 11263 185 11331 197
rect 13011 185 13079 197
rect 338 -116 409 -104
rect 338 -139 344 -116
rect 54 -198 60 -139
rect 119 -198 344 -139
rect 338 -222 344 -198
rect 403 -222 409 -116
rect 338 -234 409 -222
rect 1106 -227 1112 -175
rect 1164 -227 1170 -175
<< via1 >>
rect 13532 4884 13992 4980
rect 4129 4566 4181 4618
rect 11393 4562 11445 4614
rect 14064 4611 14116 4617
rect 14064 4571 14070 4611
rect 14070 4571 14110 4611
rect 14110 4571 14116 4611
rect 14064 4565 14116 4571
rect 14311 4660 14363 4666
rect 14311 4620 14317 4660
rect 14317 4620 14357 4660
rect 14357 4620 14363 4660
rect 14311 4614 14363 4620
rect 5126 4472 5178 4524
rect 8317 4340 9083 4436
rect 11792 4340 12558 4436
rect 5749 4244 5805 4260
rect 5749 4210 5805 4244
rect 5749 4204 5805 4210
rect 11393 4244 11445 4279
rect 11393 4227 11408 4244
rect 11408 4227 11442 4244
rect 11442 4227 11445 4244
rect 5501 4178 5553 4188
rect 5501 4136 5508 4178
rect 5508 4136 5553 4178
rect 14311 4128 14363 4180
rect 14064 4002 14116 4054
rect 6542 3796 7308 3892
rect 10037 3796 10803 3892
rect 13532 3796 13992 3892
rect 5501 3508 5553 3560
rect 14308 3558 14360 3567
rect 14308 3515 14318 3558
rect 14318 3515 14360 3558
rect 5749 3407 5805 3463
rect 14068 3479 14120 3485
rect 14068 3445 14071 3479
rect 14071 3445 14114 3479
rect 14114 3445 14120 3479
rect 14068 3433 14120 3445
rect 8317 3252 9083 3348
rect 11792 3252 12558 3348
rect 5749 3156 5805 3172
rect 5749 3122 5805 3156
rect 5749 3116 5805 3122
rect 5510 3090 5562 3100
rect 5510 3048 5556 3090
rect 5556 3048 5562 3090
rect 14308 3040 14360 3092
rect 14068 2951 14120 3003
rect 6542 2708 7308 2804
rect 10037 2708 10803 2804
rect 13532 2708 13992 2804
rect 5887 2625 5939 2677
rect 5126 2535 5178 2544
rect 5126 2501 5135 2535
rect 5135 2501 5169 2535
rect 5169 2501 5178 2535
rect 5126 2492 5178 2501
rect 4129 2461 4181 2470
rect 4129 2427 4138 2461
rect 4138 2427 4172 2461
rect 4172 2427 4181 2461
rect 4129 2418 4181 2427
rect 5250 2472 5302 2484
rect 5250 2438 5256 2472
rect 5256 2438 5296 2472
rect 5296 2438 5302 2472
rect 5250 2432 5302 2438
rect 5510 2420 5562 2472
rect 14322 2470 14374 2478
rect 14322 2426 14366 2470
rect 14366 2426 14374 2470
rect 4470 2331 4522 2383
rect 5749 2319 5805 2375
rect 14068 2391 14120 2397
rect 14068 2357 14071 2391
rect 14071 2357 14114 2391
rect 14114 2357 14120 2391
rect 14068 2345 14120 2357
rect 8317 2164 9083 2260
rect 11792 2164 12558 2260
rect 4471 2082 4523 2134
rect 5381 2084 5433 2136
rect 3725 2034 3793 2040
rect 3725 1978 3731 2034
rect 3731 1978 3787 2034
rect 3787 1978 3793 2034
rect 3725 1972 3793 1978
rect 5887 2016 5939 2068
rect 5381 1994 5433 2000
rect 5381 1954 5387 1994
rect 5387 1954 5427 1994
rect 5427 1954 5433 1994
rect 5381 1948 5433 1954
rect 14322 1952 14374 2004
rect 14068 1863 14120 1915
rect 5244 1744 5296 1796
rect 262 1620 939 1716
rect 2434 1620 3000 1716
rect 6542 1620 7308 1716
rect 10037 1620 10803 1716
rect 13532 1620 13992 1716
rect 4114 1540 4166 1592
rect 3109 1472 3161 1524
rect 4491 1540 4543 1592
rect 7976 1540 8028 1592
rect 11472 1540 11524 1592
rect 13036 1540 13088 1592
rect 15159 1540 15211 1592
rect 5872 1472 5924 1524
rect 7872 1472 7924 1524
rect 9645 1472 9697 1524
rect 11290 1472 11342 1524
rect 13223 1472 13275 1524
rect 14880 1472 14932 1524
rect 3109 1364 3161 1370
rect 3109 1324 3115 1364
rect 3115 1324 3155 1364
rect 3155 1324 3161 1364
rect 3109 1318 3161 1324
rect 4114 1382 4166 1388
rect 4114 1342 4120 1382
rect 4120 1342 4160 1382
rect 4160 1342 4166 1382
rect 4114 1333 4166 1342
rect 4491 1333 4543 1385
rect 5872 1382 5924 1388
rect 5872 1342 5878 1382
rect 5878 1342 5918 1382
rect 5918 1342 5924 1382
rect 5872 1336 5924 1342
rect 7872 1382 7924 1388
rect 7872 1342 7878 1382
rect 7878 1342 7918 1382
rect 7918 1342 7924 1382
rect 7872 1336 7924 1342
rect 7976 1382 8028 1388
rect 7976 1342 7982 1382
rect 7982 1342 8022 1382
rect 8022 1342 8028 1382
rect 7976 1336 8028 1342
rect 9645 1382 9697 1388
rect 9645 1342 9651 1382
rect 9651 1342 9691 1382
rect 9691 1342 9697 1382
rect 9645 1336 9697 1342
rect 11290 1382 11342 1388
rect 11290 1342 11296 1382
rect 11296 1342 11336 1382
rect 11336 1342 11342 1382
rect 11290 1336 11342 1342
rect 11472 1382 11524 1388
rect 11472 1342 11478 1382
rect 11478 1342 11518 1382
rect 11518 1342 11524 1382
rect 11472 1336 11524 1342
rect 13036 1382 13088 1388
rect 13036 1342 13042 1382
rect 13042 1342 13082 1382
rect 13082 1342 13088 1382
rect 13036 1336 13088 1342
rect 13223 1382 13275 1388
rect 13223 1342 13229 1382
rect 13229 1342 13269 1382
rect 13269 1342 13275 1382
rect 13223 1336 13275 1342
rect 14880 1382 14932 1388
rect 14880 1342 14886 1382
rect 14886 1342 14926 1382
rect 14926 1342 14932 1382
rect 14880 1336 14932 1342
rect 15159 1382 15211 1388
rect 15159 1342 15165 1382
rect 15165 1342 15205 1382
rect 15205 1342 15211 1382
rect 15159 1336 15211 1342
rect 3482 1295 3534 1304
rect 3482 1261 3491 1295
rect 3491 1261 3525 1295
rect 3525 1261 3534 1295
rect 3482 1252 3534 1261
rect 4679 1301 4731 1310
rect 4679 1267 4688 1301
rect 4688 1267 4722 1301
rect 4722 1267 4731 1301
rect 4679 1258 4731 1267
rect 6427 1301 6479 1310
rect 6427 1267 6436 1301
rect 6436 1267 6470 1301
rect 6470 1267 6479 1301
rect 9923 1301 9975 1310
rect 6427 1258 6479 1267
rect 8154 1287 8224 1293
rect 8154 1229 8160 1287
rect 8160 1229 8218 1287
rect 8218 1229 8224 1287
rect 8154 1223 8224 1229
rect 9923 1267 9932 1301
rect 9932 1267 9966 1301
rect 9966 1267 9975 1301
rect 9923 1258 9975 1267
rect 11650 1287 11720 1293
rect 11650 1229 11656 1287
rect 11656 1229 11714 1287
rect 11714 1229 11720 1287
rect 11650 1223 11720 1229
rect 13398 1287 13468 1293
rect 13398 1229 13404 1287
rect 13404 1229 13462 1287
rect 13462 1229 13468 1287
rect 13398 1223 13468 1229
rect 15146 1251 15198 1260
rect 15146 1217 15155 1251
rect 15155 1217 15189 1251
rect 15189 1217 15198 1251
rect 15146 1208 15198 1217
rect 1272 1076 2134 1172
rect 4798 1076 5695 1172
rect 8317 1076 9083 1172
rect 11792 1076 12558 1172
rect 2273 925 2343 931
rect 2273 867 2279 925
rect 2279 867 2337 925
rect 2337 867 2343 925
rect 2273 861 2343 867
rect 3482 916 3534 922
rect 3482 876 3488 916
rect 3488 876 3528 916
rect 3528 876 3534 916
rect 3482 870 3534 876
rect 4031 922 4083 928
rect 4031 882 4037 922
rect 4037 882 4077 922
rect 4077 882 4083 922
rect 4031 876 4083 882
rect 4679 900 4731 906
rect 4679 860 4685 900
rect 4685 860 4725 900
rect 4725 860 4731 900
rect 4679 854 4731 860
rect 5779 922 5831 928
rect 5779 882 5785 922
rect 5785 882 5825 922
rect 5825 882 5831 922
rect 5779 876 5831 882
rect 6427 900 6479 906
rect 6427 860 6433 900
rect 6433 860 6473 900
rect 6473 860 6479 900
rect 6427 854 6479 860
rect 7527 922 7579 928
rect 7527 882 7533 922
rect 7533 882 7573 922
rect 7573 882 7579 922
rect 7527 876 7579 882
rect 9275 922 9327 928
rect 9275 882 9281 922
rect 9281 882 9321 922
rect 9321 882 9327 922
rect 9275 876 9327 882
rect 8160 870 8218 876
rect 8160 824 8166 870
rect 8166 824 8212 870
rect 8212 824 8218 870
rect 8160 818 8218 824
rect 9923 900 9975 906
rect 9923 860 9929 900
rect 9929 860 9969 900
rect 9969 860 9975 900
rect 9923 854 9975 860
rect 11023 922 11075 928
rect 11023 882 11029 922
rect 11029 882 11069 922
rect 11069 882 11075 922
rect 11023 876 11075 882
rect 12771 922 12823 928
rect 12771 882 12777 922
rect 12777 882 12817 922
rect 12817 882 12823 922
rect 12771 876 12823 882
rect 14519 922 14571 928
rect 14519 882 14525 922
rect 14525 882 14565 922
rect 14565 882 14571 922
rect 14519 876 14571 882
rect 11656 870 11714 876
rect 11656 824 11662 870
rect 11662 824 11708 870
rect 11708 824 11714 870
rect 11656 818 11714 824
rect 13404 870 13462 876
rect 13404 824 13410 870
rect 13410 824 13456 870
rect 13456 824 13462 870
rect 13404 818 13462 824
rect 15146 862 15198 868
rect 15146 822 15152 862
rect 15152 822 15192 862
rect 15192 822 15198 862
rect 15146 816 15198 822
rect 3725 699 3793 767
rect 262 532 939 628
rect 2434 532 3000 628
rect 6542 532 7308 628
rect 10037 532 10803 628
rect 13532 532 13992 628
rect 60 301 119 307
rect 60 254 66 301
rect 66 254 113 301
rect 113 254 119 301
rect 60 248 119 254
rect 1112 227 1164 279
rect 2267 308 2349 314
rect 2267 238 2273 308
rect 2273 238 2343 308
rect 2343 238 2349 308
rect 2267 232 2349 238
rect 4026 311 4087 317
rect 4026 265 4032 311
rect 4032 265 4081 311
rect 4081 265 4087 311
rect 5774 311 5835 317
rect 5774 265 5780 311
rect 5780 265 5829 311
rect 5829 265 5835 311
rect 7522 311 7583 317
rect 7522 265 7528 311
rect 7528 265 7577 311
rect 7577 265 7583 311
rect 9270 311 9331 317
rect 9270 265 9276 311
rect 9276 265 9325 311
rect 9325 265 9331 311
rect 11018 311 11079 317
rect 11018 265 11024 311
rect 11024 265 11073 311
rect 11073 265 11079 311
rect 12766 311 12827 317
rect 12766 265 12772 311
rect 12772 265 12821 311
rect 12821 265 12827 311
rect 14514 311 14575 317
rect 14514 265 14520 311
rect 14520 265 14569 311
rect 14569 265 14575 311
rect 1272 -12 2134 84
rect 4798 -12 5695 84
rect 8317 -12 9083 84
rect 11792 -12 12558 84
rect 60 -198 119 -139
rect 1112 -181 1164 -175
rect 1112 -221 1118 -181
rect 1118 -221 1158 -181
rect 1158 -221 1164 -181
rect 1112 -227 1164 -221
rect 262 -556 939 -460
<< metal2 >>
rect 13532 4980 13992 4986
rect 4129 4618 4181 4624
rect 4129 4560 4181 4566
rect 11393 4614 11445 4620
rect 4138 2476 4172 4560
rect 11393 4556 11445 4562
rect 5126 4524 5178 4530
rect 5126 4466 5178 4472
rect 5135 2550 5169 4466
rect 8317 4436 9083 4442
rect 5749 4260 5805 4266
rect 5501 4188 5553 4194
rect 5501 4130 5553 4136
rect 5506 3566 5548 4130
rect 5501 3560 5553 3566
rect 5501 3502 5553 3508
rect 5749 3463 5805 4204
rect 5749 3401 5805 3407
rect 6542 3892 7308 4436
rect 5749 3172 5805 3178
rect 5510 3100 5562 3106
rect 5510 3042 5562 3048
rect 5126 2544 5178 2550
rect 5126 2486 5178 2492
rect 5250 2484 5302 2490
rect 4123 2470 4187 2476
rect 4123 2418 4129 2470
rect 4181 2418 4187 2470
rect 5515 2478 5557 3042
rect 5250 2426 5302 2432
rect 5510 2472 5562 2478
rect 4123 2412 4187 2418
rect 4470 2383 4522 2389
rect 4470 2325 4522 2331
rect 4476 2140 4517 2325
rect 4471 2134 4523 2140
rect 4471 2076 4523 2082
rect 3725 2040 3793 2046
rect 262 1716 939 1722
rect 2434 1716 3000 1722
rect 262 628 939 1081
rect 60 307 119 313
rect 60 -139 119 248
rect 60 -204 119 -198
rect 262 -460 939 532
rect 1272 1172 2134 1716
rect 1272 623 2134 1076
rect 3103 1472 3109 1524
rect 3161 1472 3167 1524
rect 3118 1376 3152 1472
rect 3109 1370 3161 1376
rect 3109 1312 3161 1318
rect 3482 1304 3534 1310
rect 3482 1246 3534 1252
rect 1112 279 1164 285
rect 1112 221 1164 227
rect 1112 -169 1163 221
rect 2273 931 2343 937
rect 2273 320 2343 861
rect 2434 628 3000 1081
rect 3491 928 3525 1246
rect 3482 922 3534 928
rect 3482 864 3534 870
rect 3491 858 3525 864
rect 3725 767 3793 1972
rect 5259 1802 5293 2426
rect 5510 2414 5562 2420
rect 5749 2375 5805 3116
rect 6542 2804 7308 3257
rect 5887 2677 5939 2683
rect 5887 2619 5939 2625
rect 5749 2313 5805 2319
rect 5381 2136 5433 2142
rect 5381 2078 5433 2084
rect 5393 2006 5421 2078
rect 5899 2068 5927 2619
rect 5881 2016 5887 2068
rect 5939 2016 5945 2068
rect 5381 2000 5433 2006
rect 5381 1942 5433 1948
rect 5244 1796 5296 1802
rect 5244 1738 5296 1744
rect 6542 1716 7308 2708
rect 4114 1592 4166 1598
rect 4114 1534 4166 1540
rect 4491 1592 4543 1598
rect 4491 1534 4543 1540
rect 4123 1394 4157 1534
rect 4114 1388 4166 1394
rect 4500 1391 4534 1534
rect 5872 1524 5924 1530
rect 5872 1466 5924 1472
rect 5881 1394 5915 1466
rect 4114 1327 4166 1333
rect 4491 1385 4543 1391
rect 4491 1327 4543 1333
rect 5872 1388 5924 1394
rect 5872 1330 5924 1336
rect 4673 1310 4737 1316
rect 4673 1258 4679 1310
rect 4731 1258 4737 1310
rect 4673 1252 4737 1258
rect 6421 1310 6485 1316
rect 6421 1258 6427 1310
rect 6479 1258 6485 1310
rect 6421 1252 6485 1258
rect 4031 928 4083 934
rect 4680 912 4730 1252
rect 4798 1172 5695 1187
rect 4031 870 4083 876
rect 4679 906 4731 912
rect 3719 699 3725 767
rect 3793 699 3799 767
rect 2261 314 2355 320
rect 2261 232 2267 314
rect 2349 232 2355 314
rect 2261 226 2355 232
rect 2434 -12 3000 532
rect 4032 317 4081 870
rect 4679 848 4731 854
rect 4798 623 5695 1076
rect 5779 928 5831 934
rect 6428 912 6478 1252
rect 8317 3348 9083 4340
rect 8317 2799 9083 3252
rect 7976 1592 8028 1598
rect 7976 1534 8028 1540
rect 7866 1472 7872 1524
rect 7924 1472 7930 1524
rect 7881 1394 7915 1472
rect 7985 1394 8019 1534
rect 7872 1388 7924 1394
rect 7872 1330 7924 1336
rect 7976 1388 8028 1394
rect 7976 1330 8028 1336
rect 8148 1293 8230 1299
rect 8148 1223 8154 1293
rect 8224 1223 8230 1293
rect 8148 1217 8230 1223
rect 5779 870 5831 876
rect 6427 906 6479 912
rect 4020 265 4026 317
rect 4087 265 4093 317
rect 5780 317 5829 870
rect 6427 848 6479 854
rect 6542 628 7308 1081
rect 7527 928 7579 934
rect 7527 870 7579 876
rect 8160 876 8218 1217
rect 5768 265 5774 317
rect 5835 265 5841 317
rect 6542 -12 7308 532
rect 7528 317 7577 870
rect 8160 812 8218 818
rect 8317 1172 9083 2164
rect 10037 3892 10803 4436
rect 11405 4279 11433 4556
rect 11792 4436 12558 4442
rect 11387 4227 11393 4279
rect 11445 4227 11451 4279
rect 10037 2804 10803 3257
rect 10037 1716 10803 2708
rect 9639 1472 9645 1524
rect 9697 1472 9703 1524
rect 9654 1394 9688 1472
rect 9645 1388 9697 1394
rect 9645 1330 9697 1336
rect 9917 1310 9981 1316
rect 9917 1258 9923 1310
rect 9975 1258 9981 1310
rect 9917 1252 9981 1258
rect 8317 623 9083 1076
rect 9275 928 9327 934
rect 9924 912 9974 1252
rect 11792 3348 12558 4340
rect 11792 2799 12558 3252
rect 11466 1540 11472 1592
rect 11524 1540 11530 1592
rect 11290 1524 11342 1530
rect 11290 1466 11342 1472
rect 11299 1394 11333 1466
rect 11481 1394 11515 1540
rect 11290 1388 11342 1394
rect 11290 1330 11342 1336
rect 11472 1388 11524 1394
rect 11472 1330 11524 1336
rect 11644 1293 11726 1299
rect 11644 1223 11650 1293
rect 11720 1223 11726 1293
rect 11644 1217 11726 1223
rect 9275 870 9327 876
rect 9923 906 9975 912
rect 7516 265 7522 317
rect 7583 265 7589 317
rect 9276 317 9325 870
rect 9923 848 9975 854
rect 10037 628 10803 1081
rect 11023 928 11075 934
rect 11023 870 11075 876
rect 11656 876 11714 1217
rect 9264 265 9270 317
rect 9331 265 9337 317
rect 10037 -12 10803 532
rect 11024 317 11073 870
rect 11656 812 11714 818
rect 11792 1172 12558 2164
rect 13532 3892 13992 4884
rect 14316 4672 14358 4705
rect 14311 4666 14363 4672
rect 14064 4617 14116 4623
rect 14311 4608 14363 4614
rect 14064 4559 14116 4565
rect 14073 4060 14107 4559
rect 14316 4186 14358 4608
rect 14311 4180 14363 4186
rect 14311 4122 14363 4128
rect 14064 4054 14116 4060
rect 14064 3996 14116 4002
rect 14308 3567 14360 3573
rect 14308 3509 14360 3515
rect 14068 3485 14120 3491
rect 14068 3427 14120 3433
rect 13532 2804 13992 3257
rect 14077 3009 14111 3427
rect 14313 3098 14355 3509
rect 14308 3092 14360 3098
rect 14308 3034 14360 3040
rect 14068 3003 14120 3009
rect 14068 2945 14120 2951
rect 13532 1716 13992 2708
rect 14322 2478 14374 2484
rect 14322 2420 14374 2426
rect 14068 2397 14120 2403
rect 14068 2339 14120 2345
rect 14077 1921 14111 2339
rect 14327 2010 14369 2420
rect 14322 2004 14374 2010
rect 14322 1946 14374 1952
rect 14068 1915 14120 1921
rect 14068 1857 14120 1863
rect 13030 1540 13036 1592
rect 13088 1540 13094 1592
rect 13045 1394 13079 1540
rect 13217 1472 13223 1524
rect 13275 1472 13281 1524
rect 13232 1394 13266 1472
rect 13036 1388 13088 1394
rect 13036 1330 13088 1336
rect 13223 1388 13275 1394
rect 13223 1330 13275 1336
rect 13392 1293 13474 1299
rect 13392 1223 13398 1293
rect 13468 1223 13474 1293
rect 13392 1217 13474 1223
rect 11792 623 12558 1076
rect 12771 928 12823 934
rect 12771 870 12823 876
rect 13404 876 13462 1217
rect 11012 265 11018 317
rect 11079 265 11085 317
rect 12772 317 12821 870
rect 13404 812 13462 818
rect 15153 1540 15159 1592
rect 15211 1540 15217 1592
rect 14874 1472 14880 1524
rect 14932 1472 14938 1524
rect 14889 1394 14923 1472
rect 15168 1394 15202 1540
rect 14880 1388 14932 1394
rect 14880 1330 14932 1336
rect 15159 1388 15211 1394
rect 15159 1330 15211 1336
rect 15140 1208 15146 1260
rect 15198 1208 15204 1260
rect 13532 628 13992 1081
rect 14519 928 14571 934
rect 14519 870 14571 876
rect 15147 874 15197 1208
rect 12760 265 12766 317
rect 12827 265 12833 317
rect 13532 -12 13992 532
rect 14520 317 14569 870
rect 15146 868 15198 874
rect 15146 810 15198 816
rect 14508 265 14514 317
rect 14575 265 14581 317
rect 1272 -18 2134 -12
rect 4798 -18 5695 -12
rect 8317 -18 9083 -12
rect 11792 -18 12558 -12
rect 1112 -175 1164 -169
rect 1112 -233 1164 -227
rect 262 -562 939 -556
<< via2 >>
rect 6542 3796 7308 3887
rect 6542 3257 7308 3796
rect 262 1620 939 1711
rect 262 1081 939 1620
rect 2434 1620 3000 1711
rect 2434 1081 3000 1620
rect 1272 84 2134 623
rect 6542 1620 7308 1711
rect 1272 -7 2134 84
rect 6542 1081 7308 1620
rect 8317 2260 9083 2799
rect 8317 2169 9083 2260
rect 4798 84 5695 623
rect 4798 -7 5695 84
rect 10037 3796 10803 3887
rect 10037 3257 10803 3796
rect 10037 1620 10803 1711
rect 10037 1081 10803 1620
rect 11792 2260 12558 2799
rect 11792 2169 12558 2260
rect 8317 84 9083 623
rect 8317 -7 9083 84
rect 13532 3796 13992 3887
rect 13532 3257 13992 3796
rect 13532 1620 13992 1711
rect 11792 84 12558 623
rect 13532 1081 13992 1620
rect 11792 -7 12558 84
<< metal3 >>
rect 5383 3887 8074 3892
rect 5383 3257 6542 3887
rect 7308 3257 8074 3887
rect 5383 3252 8074 3257
rect 14485 3252 14491 3892
rect 3727 2164 3734 2804
rect 7825 2799 14491 2804
rect 7825 2169 8317 2799
rect 9083 2169 11792 2799
rect 12558 2169 14491 2799
rect 7825 2164 14491 2169
rect 47 1711 8074 1716
rect 47 1081 262 1711
rect 939 1081 2434 1711
rect 3000 1081 6542 1711
rect 7308 1081 8074 1711
rect 47 1076 8074 1081
rect 15221 1076 15227 1716
rect 47 -12 53 628
rect 7825 623 15227 628
rect 7825 -7 8317 623
rect 9083 -7 11792 623
rect 12558 -7 15227 623
rect 7825 -12 15227 -7
<< via3 >>
rect 8074 3887 14485 3892
rect 8074 3257 10037 3887
rect 10037 3257 10803 3887
rect 10803 3257 13532 3887
rect 13532 3257 13992 3887
rect 13992 3257 14485 3887
rect 8074 3252 14485 3257
rect 3734 2164 7825 2804
rect 8074 1711 15221 1716
rect 8074 1081 10037 1711
rect 10037 1081 10803 1711
rect 10803 1081 13532 1711
rect 13532 1081 13992 1711
rect 13992 1081 15221 1711
rect 8074 1076 15221 1081
rect 53 623 7825 628
rect 53 -7 1272 623
rect 1272 -7 2134 623
rect 2134 -7 4798 623
rect 4798 -7 5695 623
rect 5695 -7 7825 623
rect 53 -12 7825 -7
<< metal4 >>
rect 47 2804 7831 4436
rect 47 2164 3734 2804
rect 7825 2164 7831 2804
rect 47 628 7831 2164
rect 47 -12 53 628
rect 7825 -12 7831 628
rect 47 -556 7831 -12
rect 8068 3892 15852 4436
rect 8068 3252 8074 3892
rect 14485 3252 15852 3892
rect 8068 1716 15852 3252
rect 8068 1076 8074 1716
rect 15221 1076 15852 1716
rect 8068 -556 15852 1076
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 28801
transform 1 0 47 0 -1 36
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 2255 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_1
timestamp 1646787781
transform -1 0 1979 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_2
timestamp 1646787781
transform -1 0 1703 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_3
timestamp 1646787781
transform -1 0 1427 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_4
timestamp 1646787781
transform -1 0 2531 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_5
timestamp 1646787781
transform -1 0 4279 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_6
timestamp 1646787781
transform -1 0 6027 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_7
timestamp 1646787781
transform -1 0 7775 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_8
timestamp 1646787781
transform -1 0 9523 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_9
timestamp 1646787781
transform -1 0 11271 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_10
timestamp 1646787781
transform -1 0 13019 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sky130_fd_sc_hd__clkbuf_1_11
timestamp 1646787781
transform -1 0 14767 0 -1 1124
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 47 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1646787781
transform 1 0 323 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1646787781
transform 1 0 599 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1646787781
transform 1 0 875 0 1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1646787781
transform -1 0 1151 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1646787781
transform -1 0 875 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1646787781
transform -1 0 599 0 -1 36
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1646787781
transform 1 0 3727 0 -1 2212
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 4003 0 -1 2212
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  sky130_fd_sc_hd__dfstp_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 5015 0 -1 2212
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 2255 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1646787781
transform 1 0 4003 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1646787781
transform 1 0 5751 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1646787781
transform 1 0 7499 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4
timestamp 1646787781
transform 1 0 9247 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_5
timestamp 1646787781
transform 1 0 10995 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_6
timestamp 1646787781
transform 1 0 12743 0 1 36
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 6947 0 -1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1646787781
transform 1 0 8419 0 -1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1646787781
transform 1 0 9983 0 -1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1646787781
transform 1 0 11455 0 -1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1646787781
transform 1 0 12927 0 -1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1646787781
transform -1 0 14399 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1646787781
transform -1 0 12927 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_8
timestamp 1646787781
transform -1 0 11455 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_9
timestamp 1646787781
transform -1 0 9891 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_10
timestamp 1646787781
transform -1 0 8419 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_11
timestamp 1646787781
transform -1 0 6947 0 1 2212
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_12
timestamp 1646787781
transform 1 0 5475 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_13
timestamp 1646787781
transform 1 0 6947 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_14
timestamp 1646787781
transform 1 0 8419 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_15
timestamp 1646787781
transform 1 0 9983 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_16
timestamp 1646787781
transform 1 0 11455 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_17
timestamp 1646787781
transform 1 0 12927 0 -1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_18
timestamp 1646787781
transform -1 0 14399 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_19
timestamp 1646787781
transform -1 0 12927 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_20
timestamp 1646787781
transform -1 0 11455 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_21
timestamp 1646787781
transform -1 0 9891 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_22
timestamp 1646787781
transform -1 0 8419 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_23
timestamp 1646787781
transform -1 0 6947 0 1 3300
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_24
timestamp 1646787781
transform 1 0 5475 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_25
timestamp 1646787781
transform 1 0 6947 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_26
timestamp 1646787781
transform 1 0 8419 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_27
timestamp 1646787781
transform 1 0 9983 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_28
timestamp 1646787781
transform 1 0 11455 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_29
timestamp 1646787781
transform 1 0 12927 0 -1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_30
timestamp 1646787781
transform -1 0 14399 0 1 4388
box -38 -48 1510 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 4739 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_1
timestamp 1646787781
transform -1 0 6487 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_2
timestamp 1646787781
transform -1 0 8235 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_3
timestamp 1646787781
transform -1 0 9983 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_4
timestamp 1646787781
transform -1 0 11731 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_5
timestamp 1646787781
transform -1 0 13479 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  sky130_fd_sc_hd__einvn_1_6
timestamp 1646787781
transform -1 0 15227 0 -1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  sky130_fd_sc_hd__einvn_4_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform -1 0 3543 0 -1 1124
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 3543 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1646787781
transform 1 0 4739 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1646787781
transform 1 0 5475 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1646787781
transform 1 0 6487 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1646787781
transform 1 0 7223 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1646787781
transform 1 0 8235 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1646787781
transform 1 0 8971 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1646787781
transform 1 0 9983 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_9
timestamp 1646787781
transform 1 0 10719 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_10
timestamp 1646787781
transform 1 0 11731 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1646787781
transform 1 0 12467 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1646787781
transform 1 0 13479 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1646787781
transform 1 0 14215 0 -1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1646787781
transform 1 0 47 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1646787781
transform 1 0 783 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1646787781
transform 1 0 1519 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1646787781
transform 1 0 2255 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_18
timestamp 1646787781
transform 1 0 2991 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_19
timestamp 1646787781
transform 1 0 3727 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_20
timestamp 1646787781
transform 1 0 4739 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_22
timestamp 1646787781
transform 1 0 6487 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_23
timestamp 1646787781
transform 1 0 7223 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_24
timestamp 1646787781
transform 1 0 8235 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_25
timestamp 1646787781
transform 1 0 8971 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_26
timestamp 1646787781
transform 1 0 9983 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_27
timestamp 1646787781
transform 1 0 10719 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_28
timestamp 1646787781
transform 1 0 11731 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_29
timestamp 1646787781
transform 1 0 12467 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_30
timestamp 1646787781
transform 1 0 13479 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_31
timestamp 1646787781
transform 1 0 14215 0 1 1124
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_32
timestamp 1646787781
transform 1 0 14491 0 1 36
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 14859 0 1 1124
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1647071613
transform 1 0 7683 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_1
timestamp 1647071613
transform 1 0 11179 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_2
timestamp 1647071613
transform 1 0 12927 0 1 1124
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  sky130_fd_sc_hd__or3_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 3083 0 1 1124
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1647018321
transform 1 0 4095 0 1 1124
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_1
timestamp 1647018321
transform 1 0 5843 0 1 1124
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_2
timestamp 1647018321
transform 1 0 9339 0 1 1124
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 1059 0 -1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1646787781
transform 1 0 1151 0 -1 36
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1646787781
transform 1 0 6487 0 -1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1646787781
transform 1 0 11731 0 -1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1646787781
transform 1 0 14215 0 -1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1646787781
transform 1 0 4923 0 -1 2212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1646787781
transform 1 0 5383 0 -1 3300
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1646787781
transform 1 0 5383 0 -1 4388
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1646787781
transform 1 0 12835 0 1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1646787781
transform 1 0 9983 0 1 1124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1646787781
transform 1 0 14399 0 1 4388
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1646787781
transform 1 0 14399 0 1 3300
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1646787781
transform 1 0 14399 0 1 2212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1646787781
transform 1 0 9891 0 1 2212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1646787781
transform 1 0 9891 0 1 3300
box -38 -48 130 592
use sky130_fd_sc_hd__xor3_1  sky130_fd_sc_hd__xor3_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 3727 0 1 2212
box -38 -48 1786 592
<< labels >>
flabel metal1 s 47 1554 76 1583 1 FreeSerif 320 0 0 0 cfg_in[0]
port 1 n
flabel metal1 s 47 1486 76 1515 1 FreeSerif 320 0 0 0 cfg_in[1]
port 2 n
flabel metal1 s 47 1418 76 1447 1 FreeSerif 320 0 0 0 cfg_in[2]
port 3 n
flabel metal1 3586 2336 3627 2377 1 FreeSerif 320 0 0 0 dout
port 4 n
flabel metal4 47 -556 7831 4436 1 FreeSerif 3200 0 0 0 GND
port 5 n
flabel metal4 8068 -556 15852 4436 1 FreeSerif 3200 0 0 0 VDD
port 6 n
flabel metal1 3587 2637 3615 2665 1 FreeSerif 320 0 0 0 n_rst
port 7 n
<< end >>
