magic
tech sky130A
magscale 1 2
timestamp 1646210680
<< nwell >>
rect -34 1604 6666 1925
<< pwell >>
rect 30 2162 74 2196
rect 766 2162 810 2196
rect 1502 2162 1546 2196
rect 2238 2162 2282 2196
rect 2974 2162 3018 2196
rect 3710 2162 3754 2196
rect 4446 2162 4490 2196
rect 5182 2162 5226 2196
rect 5918 2162 5962 2196
<< nsubdiff >>
rect 6289 1857 6323 1881
rect 6289 1773 6323 1823
rect 6289 1706 6323 1739
rect 6473 457 6507 490
rect 6473 373 6507 423
rect 6473 315 6507 339
<< nsubdiffcont >>
rect 6289 1823 6323 1857
rect 6289 1739 6323 1773
rect 6473 423 6507 457
rect 6473 339 6507 373
<< poly >>
rect 773 1494 831 1576
rect 1541 1494 1599 1576
rect 2309 1494 2367 1576
rect 4567 1420 4625 1502
<< locali >>
rect 4 2169 33 2203
rect 67 2169 125 2203
rect 159 2169 217 2203
rect 251 2169 309 2203
rect 343 2169 401 2203
rect 435 2169 493 2203
rect 527 2169 585 2203
rect 619 2169 677 2203
rect 711 2169 769 2203
rect 803 2169 861 2203
rect 895 2169 953 2203
rect 987 2169 1045 2203
rect 1079 2169 1137 2203
rect 1171 2169 1229 2203
rect 1263 2169 1321 2203
rect 1355 2169 1413 2203
rect 1447 2169 1505 2203
rect 1539 2169 1597 2203
rect 1631 2169 1689 2203
rect 1723 2169 1781 2203
rect 1815 2169 1873 2203
rect 1907 2169 1965 2203
rect 1999 2169 2057 2203
rect 2091 2169 2149 2203
rect 2183 2169 2241 2203
rect 2275 2169 2333 2203
rect 2367 2169 2425 2203
rect 2459 2169 2517 2203
rect 2551 2169 2609 2203
rect 2643 2169 2701 2203
rect 2735 2169 2793 2203
rect 2827 2169 2885 2203
rect 2919 2169 2977 2203
rect 3011 2169 3069 2203
rect 3103 2169 3161 2203
rect 3195 2169 3253 2203
rect 3287 2169 3345 2203
rect 3379 2169 3437 2203
rect 3471 2169 3529 2203
rect 3563 2169 3621 2203
rect 3655 2169 3713 2203
rect 3747 2169 3805 2203
rect 3839 2169 3897 2203
rect 3931 2169 3989 2203
rect 4023 2169 4081 2203
rect 4115 2169 4173 2203
rect 4207 2169 4265 2203
rect 4299 2169 4357 2203
rect 4391 2169 4449 2203
rect 4483 2169 4541 2203
rect 4575 2169 4633 2203
rect 4667 2169 4725 2203
rect 4759 2169 4817 2203
rect 4851 2169 4909 2203
rect 4943 2169 5001 2203
rect 5035 2169 5093 2203
rect 5127 2169 5185 2203
rect 5219 2169 5277 2203
rect 5311 2169 5369 2203
rect 5403 2169 5461 2203
rect 5495 2169 5553 2203
rect 5587 2169 5645 2203
rect 5679 2169 5737 2203
rect 5771 2169 5829 2203
rect 5863 2169 5921 2203
rect 5955 2169 6013 2203
rect 6047 2169 6105 2203
rect 6139 2169 6197 2203
rect 6231 2169 6289 2203
rect 6323 2169 6381 2203
rect 6415 2169 6473 2203
rect 6507 2169 6565 2203
rect 6599 2169 6629 2203
rect 16 1957 3260 2067
rect 3330 1957 6194 2067
rect 6277 1857 6335 1892
rect 6277 1823 6289 1857
rect 6323 1823 6335 1857
rect 6277 1773 6335 1823
rect 6277 1739 6289 1773
rect 6323 1739 6335 1773
rect 6277 1659 6335 1739
rect 6260 1625 6289 1659
rect 6323 1625 6352 1659
rect 5369 1537 6273 1591
rect 3135 1480 3823 1483
rect 3135 1424 3260 1480
rect 3330 1424 3823 1480
rect 3135 1412 3823 1424
rect 3752 1338 3823 1412
rect 5369 1338 5409 1537
rect 17 1304 3718 1329
rect 17 1264 3845 1304
rect 3594 1255 3845 1264
rect 5443 1255 5483 1454
rect 3594 1248 5483 1255
rect 3718 1164 5483 1248
rect 6461 457 6519 537
rect 6461 423 6473 457
rect 6507 423 6519 457
rect 6461 373 6519 423
rect 6461 339 6473 373
rect 6507 339 6519 373
rect 6461 304 6519 339
<< viali >>
rect 33 2169 67 2203
rect 125 2169 159 2203
rect 217 2169 251 2203
rect 309 2169 343 2203
rect 401 2169 435 2203
rect 493 2169 527 2203
rect 585 2169 619 2203
rect 677 2169 711 2203
rect 769 2169 803 2203
rect 861 2169 895 2203
rect 953 2169 987 2203
rect 1045 2169 1079 2203
rect 1137 2169 1171 2203
rect 1229 2169 1263 2203
rect 1321 2169 1355 2203
rect 1413 2169 1447 2203
rect 1505 2169 1539 2203
rect 1597 2169 1631 2203
rect 1689 2169 1723 2203
rect 1781 2169 1815 2203
rect 1873 2169 1907 2203
rect 1965 2169 1999 2203
rect 2057 2169 2091 2203
rect 2149 2169 2183 2203
rect 2241 2169 2275 2203
rect 2333 2169 2367 2203
rect 2425 2169 2459 2203
rect 2517 2169 2551 2203
rect 2609 2169 2643 2203
rect 2701 2169 2735 2203
rect 2793 2169 2827 2203
rect 2885 2169 2919 2203
rect 2977 2169 3011 2203
rect 3069 2169 3103 2203
rect 3161 2169 3195 2203
rect 3253 2169 3287 2203
rect 3345 2169 3379 2203
rect 3437 2169 3471 2203
rect 3529 2169 3563 2203
rect 3621 2169 3655 2203
rect 3713 2169 3747 2203
rect 3805 2169 3839 2203
rect 3897 2169 3931 2203
rect 3989 2169 4023 2203
rect 4081 2169 4115 2203
rect 4173 2169 4207 2203
rect 4265 2169 4299 2203
rect 4357 2169 4391 2203
rect 4449 2169 4483 2203
rect 4541 2169 4575 2203
rect 4633 2169 4667 2203
rect 4725 2169 4759 2203
rect 4817 2169 4851 2203
rect 4909 2169 4943 2203
rect 5001 2169 5035 2203
rect 5093 2169 5127 2203
rect 5185 2169 5219 2203
rect 5277 2169 5311 2203
rect 5369 2169 5403 2203
rect 5461 2169 5495 2203
rect 5553 2169 5587 2203
rect 5645 2169 5679 2203
rect 5737 2169 5771 2203
rect 5829 2169 5863 2203
rect 5921 2169 5955 2203
rect 6013 2169 6047 2203
rect 6105 2169 6139 2203
rect 6197 2169 6231 2203
rect 6289 2169 6323 2203
rect 6381 2169 6415 2203
rect 6473 2169 6507 2203
rect 6565 2169 6599 2203
rect 3260 1957 3330 2067
rect 3719 1804 3783 1872
rect 80 1724 114 1758
rect 208 1724 242 1758
rect 336 1724 370 1758
rect 464 1724 498 1758
rect 592 1724 626 1758
rect 720 1724 754 1758
rect 848 1724 882 1758
rect 976 1724 1010 1758
rect 1104 1724 1138 1758
rect 1232 1724 1266 1758
rect 1360 1724 1394 1758
rect 1488 1724 1522 1758
rect 1616 1724 1650 1758
rect 1744 1724 1778 1758
rect 1872 1724 1906 1758
rect 2000 1724 2034 1758
rect 2128 1724 2162 1758
rect 2256 1724 2290 1758
rect 2384 1724 2418 1758
rect 2512 1724 2546 1758
rect 2640 1724 2674 1758
rect 2768 1724 2802 1758
rect 2896 1724 2930 1758
rect 3024 1724 3058 1758
rect 3152 1724 3186 1758
rect 3280 1724 3314 1758
rect 3408 1724 3442 1758
rect 3536 1724 3570 1758
rect 3664 1724 3698 1758
rect 3792 1724 3826 1758
rect 3920 1724 3954 1758
rect 4048 1724 4082 1758
rect 4176 1724 4210 1758
rect 4304 1724 4338 1758
rect 4432 1724 4466 1758
rect 4560 1724 4594 1758
rect 4688 1724 4722 1758
rect 4816 1724 4850 1758
rect 4944 1724 4978 1758
rect 5072 1724 5106 1758
rect 5200 1724 5234 1758
rect 5328 1724 5362 1758
rect 5456 1724 5490 1758
rect 5584 1724 5618 1758
rect 5712 1724 5746 1758
rect 5840 1724 5874 1758
rect 5968 1724 6002 1758
rect 6096 1724 6130 1758
rect 6289 1625 6323 1659
rect 81 1526 115 1560
rect 209 1526 243 1560
rect 337 1526 371 1560
rect 465 1526 499 1560
rect 593 1526 627 1560
rect 721 1526 755 1560
rect 849 1526 883 1560
rect 977 1526 1011 1560
rect 1105 1526 1139 1560
rect 1233 1526 1267 1560
rect 1361 1526 1395 1560
rect 1489 1526 1523 1560
rect 1617 1526 1651 1560
rect 1745 1526 1779 1560
rect 1873 1526 1907 1560
rect 2001 1526 2035 1560
rect 2129 1526 2163 1560
rect 2257 1526 2291 1560
rect 2385 1526 2419 1560
rect 2513 1526 2547 1560
rect 2641 1526 2675 1560
rect 2769 1526 2803 1560
rect 2897 1526 2931 1560
rect 3025 1526 3059 1560
rect 3260 1424 3330 1480
rect 3875 1452 3909 1486
rect 4003 1452 4037 1486
rect 4131 1452 4165 1486
rect 4259 1452 4293 1486
rect 4387 1452 4421 1486
rect 4515 1452 4549 1486
rect 4643 1452 4677 1486
rect 4771 1452 4805 1486
rect 4899 1452 4933 1486
rect 5027 1452 5061 1486
rect 5155 1452 5189 1486
rect 5283 1452 5317 1486
rect 5535 1306 5569 1340
rect 5663 1306 5697 1340
rect 5791 1306 5825 1340
rect 5919 1306 5953 1340
rect 6047 1306 6081 1340
rect 6175 1306 6209 1340
rect 76 871 242 923
rect 3260 766 3330 833
rect 3260 299 3330 366
rect 76 209 242 261
<< metal1 >>
rect 4 2203 6629 2234
rect 4 2169 33 2203
rect 67 2169 125 2203
rect 159 2169 217 2203
rect 251 2169 309 2203
rect 343 2169 401 2203
rect 435 2169 493 2203
rect 527 2169 585 2203
rect 619 2169 677 2203
rect 711 2169 769 2203
rect 803 2169 861 2203
rect 895 2169 953 2203
rect 987 2169 1045 2203
rect 1079 2169 1137 2203
rect 1171 2169 1229 2203
rect 1263 2169 1321 2203
rect 1355 2169 1413 2203
rect 1447 2169 1505 2203
rect 1539 2169 1597 2203
rect 1631 2169 1689 2203
rect 1723 2169 1781 2203
rect 1815 2169 1873 2203
rect 1907 2169 1965 2203
rect 1999 2169 2057 2203
rect 2091 2169 2149 2203
rect 2183 2169 2241 2203
rect 2275 2169 2333 2203
rect 2367 2169 2425 2203
rect 2459 2169 2517 2203
rect 2551 2169 2609 2203
rect 2643 2169 2701 2203
rect 2735 2169 2793 2203
rect 2827 2169 2885 2203
rect 2919 2169 2977 2203
rect 3011 2169 3069 2203
rect 3103 2169 3161 2203
rect 3195 2169 3253 2203
rect 3287 2169 3345 2203
rect 3379 2169 3437 2203
rect 3471 2169 3529 2203
rect 3563 2169 3621 2203
rect 3655 2169 3713 2203
rect 3747 2169 3805 2203
rect 3839 2169 3897 2203
rect 3931 2169 3989 2203
rect 4023 2169 4081 2203
rect 4115 2169 4173 2203
rect 4207 2169 4265 2203
rect 4299 2169 4357 2203
rect 4391 2169 4449 2203
rect 4483 2169 4541 2203
rect 4575 2169 4633 2203
rect 4667 2169 4725 2203
rect 4759 2169 4817 2203
rect 4851 2169 4909 2203
rect 4943 2169 5001 2203
rect 5035 2169 5093 2203
rect 5127 2169 5185 2203
rect 5219 2169 5277 2203
rect 5311 2169 5369 2203
rect 5403 2169 5461 2203
rect 5495 2169 5553 2203
rect 5587 2169 5645 2203
rect 5679 2169 5737 2203
rect 5771 2169 5829 2203
rect 5863 2169 5921 2203
rect 5955 2169 6013 2203
rect 6047 2169 6105 2203
rect 6139 2169 6197 2203
rect 6231 2169 6289 2203
rect 6323 2169 6381 2203
rect 6415 2169 6473 2203
rect 6507 2169 6565 2203
rect 6599 2169 6629 2203
rect 4 2138 6629 2169
rect 3254 2067 3336 2079
rect 3250 1957 3260 2067
rect 3330 1957 3340 2067
rect 3254 1945 3336 1957
rect 3713 1872 3789 1884
rect 3709 1801 3719 1872
rect 3783 1801 3793 1872
rect 3713 1792 3789 1801
rect 4 1758 6628 1764
rect 4 1724 80 1758
rect 114 1724 208 1758
rect 242 1724 336 1758
rect 370 1724 464 1758
rect 498 1724 592 1758
rect 626 1724 720 1758
rect 754 1724 848 1758
rect 882 1724 976 1758
rect 1010 1724 1104 1758
rect 1138 1724 1232 1758
rect 1266 1724 1360 1758
rect 1394 1724 1488 1758
rect 1522 1724 1616 1758
rect 1650 1724 1744 1758
rect 1778 1724 1872 1758
rect 1906 1724 2000 1758
rect 2034 1724 2128 1758
rect 2162 1724 2256 1758
rect 2290 1724 2384 1758
rect 2418 1724 2512 1758
rect 2546 1724 2640 1758
rect 2674 1724 2768 1758
rect 2802 1724 2896 1758
rect 2930 1724 3024 1758
rect 3058 1724 3152 1758
rect 3186 1724 3280 1758
rect 3314 1724 3408 1758
rect 3442 1724 3536 1758
rect 3570 1724 3664 1758
rect 3698 1724 3792 1758
rect 3826 1724 3920 1758
rect 3954 1724 4048 1758
rect 4082 1724 4176 1758
rect 4210 1724 4304 1758
rect 4338 1724 4432 1758
rect 4466 1724 4560 1758
rect 4594 1724 4688 1758
rect 4722 1724 4816 1758
rect 4850 1724 4944 1758
rect 4978 1724 5072 1758
rect 5106 1724 5200 1758
rect 5234 1724 5328 1758
rect 5362 1724 5456 1758
rect 5490 1724 5584 1758
rect 5618 1724 5712 1758
rect 5746 1724 5840 1758
rect 5874 1724 5968 1758
rect 6002 1724 6096 1758
rect 6130 1724 6628 1758
rect 4 1718 6628 1724
rect 6260 1659 6352 1690
rect 6260 1625 6289 1659
rect 6323 1625 6352 1659
rect 6260 1594 6352 1625
rect 4 1560 6628 1566
rect 4 1526 81 1560
rect 115 1526 209 1560
rect 243 1526 337 1560
rect 371 1526 465 1560
rect 499 1526 593 1560
rect 627 1526 721 1560
rect 755 1526 849 1560
rect 883 1526 977 1560
rect 1011 1526 1105 1560
rect 1139 1526 1233 1560
rect 1267 1526 1361 1560
rect 1395 1526 1489 1560
rect 1523 1526 1617 1560
rect 1651 1526 1745 1560
rect 1779 1526 1873 1560
rect 1907 1526 2001 1560
rect 2035 1526 2129 1560
rect 2163 1526 2257 1560
rect 2291 1526 2385 1560
rect 2419 1526 2513 1560
rect 2547 1526 2641 1560
rect 2675 1526 2769 1560
rect 2803 1526 2897 1560
rect 2931 1526 3025 1560
rect 3059 1526 6628 1560
rect 4 1520 6628 1526
rect 3254 1480 3336 1492
rect 3254 1412 3260 1480
rect 3330 1412 3336 1480
rect 3364 1486 6318 1492
rect 3364 1452 3875 1486
rect 3909 1452 4003 1486
rect 4037 1452 4131 1486
rect 4165 1452 4259 1486
rect 4293 1452 4387 1486
rect 4421 1452 4515 1486
rect 4549 1452 4643 1486
rect 4677 1452 4771 1486
rect 4805 1452 4899 1486
rect 4933 1452 5027 1486
rect 5061 1452 5155 1486
rect 5189 1452 5283 1486
rect 5317 1452 6318 1486
rect 3364 1446 6318 1452
rect 3364 1384 3410 1446
rect 4 1338 3410 1384
rect 6272 1384 6318 1446
rect 3471 1340 6227 1346
rect 3471 1310 5535 1340
rect 4 1306 5535 1310
rect 5569 1306 5663 1340
rect 5697 1306 5791 1340
rect 5825 1306 5919 1340
rect 5953 1306 6047 1340
rect 6081 1306 6175 1340
rect 6209 1310 6227 1340
rect 6272 1338 6628 1384
rect 6209 1306 6628 1310
rect 4 1300 6628 1306
rect 4 1264 3517 1300
rect 3700 1249 3783 1270
rect 6181 1264 6628 1300
rect 3700 1230 3719 1249
rect 3256 1174 3266 1230
rect 3330 1174 3340 1230
rect 3709 1193 3719 1230
rect 3752 1174 3783 1193
rect 2 923 254 929
rect 2 871 76 923
rect 242 871 254 923
rect 2 865 254 871
rect 3248 833 3342 839
rect 3248 766 3260 833
rect 3330 766 3342 833
rect 3248 760 3342 766
rect 6536 571 6628 602
rect 6536 537 6565 571
rect 6599 537 6628 571
rect 6536 506 6628 537
rect 3248 366 3342 372
rect 3248 299 3260 366
rect 3330 299 3342 366
rect 3248 293 3342 299
rect 64 261 254 267
rect 64 209 76 261
rect 242 209 254 261
rect 64 203 254 209
<< via1 >>
rect 3260 1957 3330 2067
rect 3719 1804 3783 1872
rect 3719 1801 3783 1804
rect 3260 1424 3330 1480
rect 3260 1412 3330 1424
rect 3266 1174 3330 1230
rect 3719 1193 3783 1249
rect 76 871 242 923
rect 3260 766 3330 833
rect 3260 299 3330 366
rect 76 209 242 261
<< metal2 >>
rect 3260 2067 3330 2073
rect 3260 1480 3330 1957
rect 3260 1230 3330 1412
rect 3260 1174 3266 1230
rect 3719 1872 3783 1882
rect 3719 1249 3783 1801
rect 3719 1183 3783 1193
rect 76 923 242 933
rect 76 261 242 871
rect 3260 833 3330 1174
rect 3260 366 3330 766
rect 3260 289 3330 299
rect 76 199 242 209
use p-leg_fet_16  p-leg_fet_16_4 ~/proj/sstl-design/layout
timestamp 1643664681
transform 1 0 3103 0 -1 769
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_1
timestamp 1643664681
transform 1 0 3103 0 1 363
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_3
timestamp 1643664681
transform 1 0 1055 0 -1 769
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_0
timestamp 1643664681
transform 1 0 1055 0 1 363
box -1089 -161 1089 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 4 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1644111581
transform 1 0 740 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1644111581
transform 1 0 1476 0 1 10
box -38 -48 774 592
use p-leg_fet_16  p-leg_fet_16_5
timestamp 1643664681
transform 1 0 5151 0 -1 769
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_2
timestamp 1643664681
transform 1 0 5151 0 1 363
box -1089 -161 1089 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1644111581
transform 1 0 2212 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1644111581
transform 1 0 2948 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1644111581
transform 1 0 3684 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1644111581
transform 1 0 4420 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1644111581
transform 1 0 5156 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1644111581
transform 1 0 5892 0 1 10
box -38 -48 774 592
use p-leg_6  p-leg_6_2 ~/proj/sstl-design/layout
timestamp 1643158822
transform 1 0 2594 0 -1 1415
box -1089 -161 -191 198
use p-leg_6  p-leg_6_1
timestamp 1643158822
transform 1 0 1826 0 -1 1415
box -1089 -161 -191 198
use p-leg_6  p-leg_6_0
timestamp 1643158822
transform 1 0 1058 0 -1 1415
box -1089 -161 -191 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_10
timestamp 1644111581
transform 1 0 740 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_9
timestamp 1644111581
transform 1 0 4 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1644111581
transform 1 0 1476 0 1 1098
box -38 -48 774 592
use p-leg_polyres  p-leg_polyres_0 ~/proj/sstl-design/layout
timestamp 1643152784
transform 0 -1 3515 1 0 1197
box -33 -253 33 253
use p-leg_6  p-leg_6_4
timestamp 1643158822
transform 1 0 4852 0 -1 1341
box -1089 -161 -191 198
use p-leg_6  p-leg_6_3
timestamp 1643158822
transform 1 0 3362 0 -1 1415
box -1089 -161 -191 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1644111581
transform 1 0 2948 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1644111581
transform 1 0 2212 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1644111581
transform 1 0 3684 0 1 1098
box -38 -48 774 592
use p-leg_6  p-leg_6_5
timestamp 1643158822
transform 1 0 5620 0 -1 1341
box -1089 -161 -191 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1644111581
transform 1 0 5156 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1644111581
transform 1 0 4420 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1644111581
transform 1 0 5892 0 1 1098
box -38 -48 774 592
use p-leg_fet_16  p-leg_fet_16_8
timestamp 1643664681
transform -1 0 1057 0 1 1869
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_6
timestamp 1643664681
transform -1 0 3105 0 1 1869
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_7
timestamp 1643664681
transform -1 0 5153 0 1 1869
box -1089 -161 1089 198
use p-leg_6  p-leg_6_6
timestamp 1643158822
transform 1 0 6512 0 1 1451
box -1089 -161 -191 198
<< labels >>
flabel metal1 s 30 553 30 553 7 FreeSerif 640 0 0 0 VDD
port 3 w
flabel metal1 s 30 1641 30 1641 7 FreeSerif 640 0 0 0 VDD
port 3 w
flabel metal1 s 26 1740 26 1740 7 FreeSerif 640 0 0 0 n_cal_ctrl[0]
port 4 w
flabel metal1 s 27 1542 27 1542 7 FreeSerif 640 0 0 0 n_cal_ctrl[1]
port 5 w
flabel metal1 3294 997 3294 997 7 FreeSerif 640 0 0 0 v_pullup
flabel metal2 s 3752 1250 3752 1250 3 FreeSerif 640 0 0 0 DQ
port 2 e
flabel metal1 s 27 1286 27 1286 7 FreeSerif 640 0 0 0 n_cal_ctrl[3]
port 7 w
flabel metal1 s 27 1360 27 1360 7 FreeSerif 640 0 0 0 n_cal_ctrl[2]
port 6 w
flabel metal1 s 2 865 2 929 7 FreeSerif 800 0 0 0 n_pu_ctrl
port 8 w
<< end >>
