magic
tech sky130A
magscale 1 2
timestamp 1646794558
<< checkpaint >>
rect 11573 647465 53167 689591
rect 3138 647230 58204 647465
rect 3068 638726 58296 647230
rect 3138 638579 58204 638726
<< metal1 >>
rect 7241 643202 7251 643298
rect 7469 643202 7479 643298
rect 8713 643202 8723 643298
rect 8941 643202 8951 643298
rect 10185 643202 10195 643298
rect 10413 643202 10423 643298
rect 11657 643202 11667 643298
rect 11885 643202 11895 643298
rect 13129 643202 13139 643298
rect 13357 643202 13367 643298
rect 14601 643202 14611 643298
rect 14829 643202 14839 643298
rect 16073 643202 16083 643298
rect 16301 643202 16311 643298
rect 17545 643202 17555 643298
rect 17773 643202 17783 643298
rect 19017 643202 19027 643298
rect 19245 643202 19255 643298
rect 20489 643202 20499 643298
rect 20717 643202 20727 643298
rect 21961 643202 21971 643298
rect 22189 643202 22199 643298
rect 23433 643202 23443 643298
rect 23661 643202 23671 643298
rect 24905 643202 24915 643298
rect 25133 643202 25143 643298
rect 26377 643202 26387 643298
rect 26605 643202 26615 643298
rect 27849 643202 27859 643298
rect 28077 643202 28087 643298
rect 29321 643202 29331 643298
rect 29549 643202 29559 643298
rect 30793 643202 30803 643298
rect 31021 643202 31031 643298
rect 32265 643202 32275 643298
rect 32493 643202 32503 643298
rect 33737 643202 33747 643298
rect 33965 643202 33975 643298
rect 35209 643202 35219 643298
rect 35437 643202 35447 643298
rect 36681 643202 36691 643298
rect 36909 643202 36919 643298
rect 38153 643202 38163 643298
rect 38381 643202 38391 643298
rect 39625 643202 39635 643298
rect 39853 643202 39863 643298
rect 41097 643202 41107 643298
rect 41325 643202 41335 643298
rect 42569 643202 42579 643298
rect 42797 643202 42807 643298
rect 44041 643202 44051 643298
rect 44269 643202 44279 643298
rect 45513 643202 45523 643298
rect 45741 643202 45751 643298
rect 46985 643202 46995 643298
rect 47213 643202 47223 643298
rect 48457 643202 48467 643298
rect 48685 643202 48695 643298
rect 49929 643202 49939 643298
rect 50157 643202 50167 643298
rect 51401 643202 51411 643298
rect 51629 643202 51639 643298
rect 52873 643202 52883 643298
rect 53101 643202 53111 643298
rect 54315 642961 57514 643052
rect 54228 642917 57514 642961
rect 54315 642827 57514 642917
rect 57739 642827 57745 643052
rect 7241 642658 7251 642754
rect 7469 642658 7479 642754
rect 8713 642658 8723 642754
rect 8941 642658 8951 642754
rect 10185 642658 10195 642754
rect 10413 642658 10423 642754
rect 11657 642658 11667 642754
rect 11885 642658 11895 642754
rect 13129 642658 13139 642754
rect 13357 642658 13367 642754
rect 14601 642658 14611 642754
rect 14829 642658 14839 642754
rect 16073 642658 16083 642754
rect 16301 642658 16311 642754
rect 17545 642658 17555 642754
rect 17773 642658 17783 642754
rect 19017 642658 19027 642754
rect 19245 642658 19255 642754
rect 20489 642658 20499 642754
rect 20717 642658 20727 642754
rect 21961 642658 21971 642754
rect 22189 642658 22199 642754
rect 23433 642658 23443 642754
rect 23661 642658 23671 642754
rect 24905 642658 24915 642754
rect 25133 642658 25143 642754
rect 26377 642658 26387 642754
rect 26605 642658 26615 642754
rect 27849 642658 27859 642754
rect 28077 642658 28087 642754
rect 29321 642658 29331 642754
rect 29549 642658 29559 642754
rect 30793 642658 30803 642754
rect 31021 642658 31031 642754
rect 32265 642658 32275 642754
rect 32493 642658 32503 642754
rect 33737 642658 33747 642754
rect 33965 642658 33975 642754
rect 35209 642658 35219 642754
rect 35437 642658 35447 642754
rect 36681 642658 36691 642754
rect 36909 642658 36919 642754
rect 38153 642658 38163 642754
rect 38381 642658 38391 642754
rect 39625 642658 39635 642754
rect 39853 642658 39863 642754
rect 41097 642658 41107 642754
rect 41325 642658 41335 642754
rect 42569 642658 42579 642754
rect 42797 642658 42807 642754
rect 44041 642658 44051 642754
rect 44269 642658 44279 642754
rect 45513 642658 45523 642754
rect 45741 642658 45751 642754
rect 46985 642658 46995 642754
rect 47213 642658 47223 642754
rect 48457 642658 48467 642754
rect 48685 642658 48695 642754
rect 49929 642658 49939 642754
rect 50157 642658 50167 642754
rect 51401 642658 51411 642754
rect 51629 642658 51639 642754
rect 52873 642658 52883 642754
rect 53101 642658 53111 642754
<< via1 >>
rect 7251 643202 7469 643298
rect 8723 643202 8941 643298
rect 10195 643202 10413 643298
rect 11667 643202 11885 643298
rect 13139 643202 13357 643298
rect 14611 643202 14829 643298
rect 16083 643202 16301 643298
rect 17555 643202 17773 643298
rect 19027 643202 19245 643298
rect 20499 643202 20717 643298
rect 21971 643202 22189 643298
rect 23443 643202 23661 643298
rect 24915 643202 25133 643298
rect 26387 643202 26605 643298
rect 27859 643202 28077 643298
rect 29331 643202 29549 643298
rect 30803 643202 31021 643298
rect 32275 643202 32493 643298
rect 33747 643202 33965 643298
rect 35219 643202 35437 643298
rect 36691 643202 36909 643298
rect 38163 643202 38381 643298
rect 39635 643202 39853 643298
rect 41107 643202 41325 643298
rect 42579 643202 42797 643298
rect 44051 643202 44269 643298
rect 45523 643202 45741 643298
rect 46995 643202 47213 643298
rect 48467 643202 48685 643298
rect 49939 643202 50157 643298
rect 51411 643202 51629 643298
rect 52883 643202 53101 643298
rect 57514 642827 57739 643052
rect 7251 642658 7469 642754
rect 8723 642658 8941 642754
rect 10195 642658 10413 642754
rect 11667 642658 11885 642754
rect 13139 642658 13357 642754
rect 14611 642658 14829 642754
rect 16083 642658 16301 642754
rect 17555 642658 17773 642754
rect 19027 642658 19245 642754
rect 20499 642658 20717 642754
rect 21971 642658 22189 642754
rect 23443 642658 23661 642754
rect 24915 642658 25133 642754
rect 26387 642658 26605 642754
rect 27859 642658 28077 642754
rect 29331 642658 29549 642754
rect 30803 642658 31021 642754
rect 32275 642658 32493 642754
rect 33747 642658 33965 642754
rect 35219 642658 35437 642754
rect 36691 642658 36909 642754
rect 38163 642658 38381 642754
rect 39635 642658 39853 642754
rect 41107 642658 41325 642754
rect 42579 642658 42797 642754
rect 44051 642658 44269 642754
rect 45523 642658 45741 642754
rect 46995 642658 47213 642754
rect 48467 642658 48685 642754
rect 49939 642658 50157 642754
rect 51411 642658 51629 642754
rect 52883 642658 53101 642754
<< metal2 >>
rect 45991 687785 46650 687794
rect 31964 687750 32623 687759
rect 31964 680231 32623 687091
rect 45991 679877 46650 687126
rect 201295 675703 201384 675805
rect 215296 675654 215385 675823
rect 14344 669979 14353 670638
rect 15012 669979 22362 670638
rect 21703 667744 22362 669979
rect 15653 645391 15712 645799
rect 8492 645332 15712 645391
rect 7251 643298 7469 643308
rect 8554 643242 8594 645332
rect 15773 645244 15832 645876
rect 9918 645185 15832 645244
rect 8723 643298 8941 643308
rect 7251 643192 7469 643202
rect 10026 643237 10066 645185
rect 15893 645086 15952 645599
rect 11315 645027 15952 645086
rect 10195 643298 10413 643308
rect 8723 643192 8941 643202
rect 11498 643242 11538 645027
rect 12970 644927 13010 644933
rect 16013 644927 16072 645797
rect 12968 644868 16072 644927
rect 11667 643298 11885 643308
rect 10195 643192 10413 643202
rect 12970 643247 13010 644868
rect 16133 644745 16192 645679
rect 14386 644686 16192 644745
rect 13139 643298 13357 643308
rect 11667 643192 11885 643202
rect 14442 643258 14482 644686
rect 16253 644536 16312 645609
rect 15904 644477 16312 644536
rect 16373 644546 16432 645724
rect 16373 644487 17455 644546
rect 14611 643298 14829 643308
rect 13139 643192 13357 643202
rect 15914 643232 15954 644477
rect 16083 643298 16301 643308
rect 14611 643192 14829 643202
rect 17386 643222 17426 644487
rect 18529 643461 18587 645573
rect 18805 643602 18863 645588
rect 19080 643727 19138 645568
rect 19355 643847 19413 645578
rect 19912 643992 19970 645593
rect 20032 644087 20090 645688
rect 20152 644202 20210 645648
rect 20272 644302 20330 645578
rect 26143 645289 26429 645293
rect 26555 645289 26629 645582
rect 26138 645284 26629 645289
rect 26138 644998 26143 645284
rect 26429 644998 26629 645284
rect 26138 644993 26629 644998
rect 26143 644989 26429 644993
rect 26555 644971 26629 644993
rect 26670 644853 26702 645540
rect 26740 645324 26789 645557
rect 26740 645226 26937 645324
rect 26789 645146 26937 645226
rect 26789 644989 26937 644998
rect 26349 644819 26702 644853
rect 26349 644696 26370 644819
rect 26350 644507 26370 644635
rect 26682 644507 26702 644819
rect 26350 644490 26702 644507
rect 26670 644481 26702 644490
rect 27034 644499 27094 645568
rect 27592 644600 27652 645600
rect 33996 645431 34054 645576
rect 33577 645373 34054 645431
rect 27592 644540 32250 644600
rect 27034 644439 30707 644499
rect 20272 644244 29228 644302
rect 20152 644144 27767 644202
rect 20032 644029 26341 644087
rect 19912 643934 24831 643992
rect 19355 643789 23350 643847
rect 19080 643669 21879 643727
rect 18805 643544 20398 643602
rect 18529 643403 18977 643461
rect 17555 643298 17773 643308
rect 16083 643192 16301 643202
rect 18858 643229 18898 643403
rect 19027 643298 19245 643308
rect 17555 643192 17773 643202
rect 20330 643245 20370 643544
rect 20499 643298 20717 643308
rect 19027 643192 19245 643202
rect 21802 643241 21842 643669
rect 21971 643298 22189 643308
rect 20499 643192 20717 643202
rect 23274 643231 23314 643789
rect 23443 643298 23661 643308
rect 21971 643192 22189 643202
rect 24746 643236 24786 643934
rect 24915 643298 25133 643308
rect 23443 643192 23661 643202
rect 26218 643236 26258 644029
rect 26387 643298 26605 643308
rect 24915 643192 25133 643202
rect 27690 643236 27730 644144
rect 27859 643298 28077 643308
rect 26387 643192 26605 643202
rect 29162 643236 29202 644244
rect 29331 643298 29549 643308
rect 27859 643192 28077 643202
rect 30634 643241 30674 644439
rect 30803 643298 31021 643308
rect 29331 643192 29549 643202
rect 32106 643252 32146 644540
rect 32275 643298 32493 643308
rect 30803 643192 31021 643202
rect 33578 643225 33618 645373
rect 34116 643470 34174 645566
rect 34236 643593 34294 645593
rect 34356 643715 34414 645566
rect 34913 643844 34971 645566
rect 35188 643961 35246 645582
rect 35463 644090 35521 645582
rect 35739 644196 35797 645582
rect 38453 644322 38509 645575
rect 38545 644458 38601 645564
rect 38637 644572 38693 645575
rect 38729 644709 38785 645575
rect 38821 644823 38877 645575
rect 38913 644914 38969 645586
rect 39005 645017 39061 645564
rect 39005 644961 54301 645017
rect 38913 644858 52979 644914
rect 38821 644767 51282 644823
rect 38729 644653 49903 644709
rect 38637 644516 48365 644572
rect 38545 644402 46919 644458
rect 38453 644321 45378 644322
rect 38453 644266 45394 644321
rect 35739 644138 43929 644196
rect 35463 644032 42499 644090
rect 35188 643903 41012 643961
rect 34913 643786 39537 643844
rect 34356 643657 38045 643715
rect 34236 643535 36636 643593
rect 34116 643412 35150 643470
rect 33747 643298 33965 643308
rect 32275 643192 32493 643202
rect 33747 643192 33965 643202
rect 35050 643162 35090 643412
rect 35219 643298 35437 643308
rect 35219 643192 35437 643202
rect 36522 643105 36562 643535
rect 36691 643298 36909 643308
rect 36691 643192 36909 643202
rect 37994 643100 38034 643657
rect 38163 643298 38381 643308
rect 38163 643192 38381 643202
rect 39466 643088 39506 643786
rect 39635 643298 39853 643308
rect 39635 643192 39853 643202
rect 40938 643026 40978 643903
rect 41107 643298 41325 643308
rect 42410 643230 42450 644032
rect 42579 643298 42797 643308
rect 41107 643192 41325 643202
rect 42579 643192 42797 643202
rect 43882 643196 43922 644138
rect 44051 643298 44269 643308
rect 44051 643192 44269 643202
rect 45354 643146 45394 644266
rect 45523 643298 45741 643308
rect 45523 643192 45741 643202
rect 46826 643129 46866 644402
rect 46995 643298 47213 643308
rect 46995 643192 47213 643202
rect 48298 643137 48338 644516
rect 48467 643298 48685 643308
rect 48467 643192 48685 643202
rect 49770 643096 49810 644653
rect 49939 643298 50157 643308
rect 49939 643192 50157 643202
rect 51242 643120 51282 644767
rect 51411 643298 51629 643308
rect 51411 643192 51629 643202
rect 52714 643021 52754 644858
rect 52883 643298 53101 643308
rect 52883 643192 53101 643202
rect 54186 643102 54226 644961
rect 57514 643052 57739 643069
rect 7251 642754 7469 642764
rect 7082 642601 7122 642699
rect 7251 642648 7469 642658
rect 8723 642754 8941 642764
rect 8723 642648 8941 642658
rect 10195 642754 10413 642764
rect 10195 642648 10413 642658
rect 11667 642754 11885 642764
rect 11667 642648 11885 642658
rect 13139 642754 13357 642764
rect 13139 642648 13357 642658
rect 14611 642754 14829 642764
rect 14611 642648 14829 642658
rect 16083 642754 16301 642764
rect 16083 642648 16301 642658
rect 17555 642754 17773 642764
rect 17555 642648 17773 642658
rect 19027 642754 19245 642764
rect 19027 642648 19245 642658
rect 20499 642754 20717 642764
rect 20499 642648 20717 642658
rect 21971 642754 22189 642764
rect 21971 642648 22189 642658
rect 23443 642754 23661 642764
rect 23443 642648 23661 642658
rect 24915 642754 25133 642764
rect 24915 642648 25133 642658
rect 26387 642754 26605 642764
rect 26387 642648 26605 642658
rect 27859 642754 28077 642764
rect 27859 642648 28077 642658
rect 29331 642754 29549 642764
rect 29331 642648 29549 642658
rect 30803 642754 31021 642764
rect 30803 642648 31021 642658
rect 32275 642754 32493 642764
rect 32275 642648 32493 642658
rect 33747 642754 33965 642764
rect 33747 642648 33965 642658
rect 35219 642754 35437 642764
rect 35219 642648 35437 642658
rect 36691 642754 36909 642764
rect 36691 642648 36909 642658
rect 38163 642754 38381 642764
rect 38163 642648 38381 642658
rect 39635 642754 39853 642764
rect 39635 642648 39853 642658
rect 41107 642754 41325 642764
rect 41107 642648 41325 642658
rect 42579 642754 42797 642764
rect 42579 642648 42797 642658
rect 44051 642754 44269 642764
rect 44051 642648 44269 642658
rect 45523 642754 45741 642764
rect 45523 642648 45741 642658
rect 46995 642754 47213 642764
rect 46995 642648 47213 642658
rect 48467 642754 48685 642764
rect 48467 642648 48685 642658
rect 49939 642754 50157 642764
rect 49939 642648 50157 642658
rect 51411 642754 51629 642764
rect 51411 642648 51629 642658
rect 52883 642754 53101 642764
rect 52883 642648 53101 642658
rect 6999 641447 7206 642601
rect 57514 641802 57739 642827
rect 57514 641568 57739 641577
rect 6999 641231 7206 641240
rect 126679 3554 127384 4191
rect 126679 3530 127435 3554
rect 126679 2835 126731 3530
rect 127426 2835 127435 3530
rect 126679 2820 127435 2835
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 213
rect 126679 6 127384 2820
rect 126998 -800 127110 6
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 31964 687091 32623 687750
rect 45991 687126 46650 687785
rect 14353 669979 15012 670638
rect 7251 643202 7469 643298
rect 8723 643202 8941 643298
rect 10195 643202 10413 643298
rect 11667 643202 11885 643298
rect 13139 643202 13357 643298
rect 14611 643202 14829 643298
rect 16083 643202 16301 643298
rect 26143 644998 26429 645284
rect 26789 644998 26937 645146
rect 26370 644507 26682 644819
rect 17555 643202 17773 643298
rect 19027 643202 19245 643298
rect 20499 643202 20717 643298
rect 21971 643202 22189 643298
rect 23443 643202 23661 643298
rect 24915 643202 25133 643298
rect 26387 643202 26605 643298
rect 27859 643202 28077 643298
rect 29331 643202 29549 643298
rect 30803 643202 31021 643298
rect 32275 643202 32493 643298
rect 33747 643202 33965 643298
rect 35219 643202 35437 643298
rect 36691 643202 36909 643298
rect 38163 643202 38381 643298
rect 39635 643202 39853 643298
rect 41107 643202 41325 643298
rect 42579 643202 42797 643298
rect 44051 643202 44269 643298
rect 45523 643202 45741 643298
rect 46995 643202 47213 643298
rect 48467 643202 48685 643298
rect 49939 643202 50157 643298
rect 51411 643202 51629 643298
rect 52883 643202 53101 643298
rect 7251 642658 7469 642754
rect 8723 642658 8941 642754
rect 10195 642658 10413 642754
rect 11667 642658 11885 642754
rect 13139 642658 13357 642754
rect 14611 642658 14829 642754
rect 16083 642658 16301 642754
rect 17555 642658 17773 642754
rect 19027 642658 19245 642754
rect 20499 642658 20717 642754
rect 21971 642658 22189 642754
rect 23443 642658 23661 642754
rect 24915 642658 25133 642754
rect 26387 642658 26605 642754
rect 27859 642658 28077 642754
rect 29331 642658 29549 642754
rect 30803 642658 31021 642754
rect 32275 642658 32493 642754
rect 33747 642658 33965 642754
rect 35219 642658 35437 642754
rect 36691 642658 36909 642754
rect 38163 642658 38381 642754
rect 39635 642658 39853 642754
rect 41107 642658 41325 642754
rect 42579 642658 42797 642754
rect 44051 642658 44269 642754
rect 45523 642658 45741 642754
rect 46995 642658 47213 642754
rect 48467 642658 48685 642754
rect 49939 642658 50157 642754
rect 51411 642658 51629 642754
rect 52883 642658 53101 642754
rect 57514 641577 57739 641802
rect 6999 641240 7206 641447
rect 126731 2835 127426 3530
<< metal3 >>
rect 16194 702300 21194 704800
rect 18694 688664 21194 702300
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 68194 688671 70694 702300
rect 165676 701964 170594 702300
rect 170894 701964 173094 704800
rect 173394 702477 175594 704800
rect 165676 699764 173094 701964
rect 165676 693758 170594 699764
rect 173298 699486 175798 702477
rect 173298 696988 173299 699486
rect 175797 696988 175798 699486
rect 173298 696865 175798 696988
rect 175894 693758 180894 704800
rect 217294 699492 222294 704800
rect 222594 703413 224794 704800
rect 222482 702159 224982 703413
rect 222477 699661 222483 702159
rect 224981 699661 224987 702159
rect 225094 701830 227294 704800
rect 227594 704448 232594 704800
rect 227594 702300 232595 704448
rect 227663 701830 232595 702300
rect 222482 699660 224982 699661
rect 225094 699630 232595 701830
rect 217176 699487 222294 699492
rect 227663 699487 232595 699630
rect 318994 699585 323994 704800
rect 324294 702094 326494 704800
rect 326794 702122 328994 704800
rect 329294 702122 334294 704800
rect 326794 699922 334294 702122
rect 324294 699888 326494 699894
rect 329294 699585 334294 699922
rect 217176 699486 232595 699487
rect 219674 696990 232595 699486
rect 318700 697085 334294 699585
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 413394 702099 415894 702300
rect 413394 702093 416035 702099
rect 413394 699895 413837 702093
rect 413394 699889 416035 699895
rect 217176 696982 219674 696988
rect 219794 696987 232595 696990
rect 164546 691258 172231 693758
rect 174731 691258 180894 693758
rect 178394 691256 180894 691258
rect 18694 687750 33489 688664
rect 18694 687091 31964 687750
rect 32623 687091 33489 687750
rect 18694 686164 33489 687091
rect 44999 687785 70694 688671
rect 44999 687126 45991 687785
rect 46650 687126 70694 687785
rect 44999 686171 70694 687126
rect 18694 686083 21194 686164
rect -800 682742 1700 685242
rect -800 680242 12279 682742
rect 9779 671807 12279 680242
rect 9779 670638 15560 671807
rect 9779 669979 14353 670638
rect 15012 669979 15560 670638
rect 9779 669307 15560 669979
rect 326068 657980 328568 697085
rect 329294 697047 331794 697085
rect 49676 656363 331553 657980
rect 48111 655930 49833 656363
rect 50266 655930 331553 656363
rect 49676 655928 331553 655930
rect 413394 655832 415894 699889
rect 582300 677984 584800 682984
rect 47359 655405 419024 655832
rect 49671 654203 419024 655405
rect 49671 653776 50443 654203
rect 50870 653776 419024 654203
rect 49671 653743 419024 653776
rect -800 643842 1660 648642
rect 24904 645288 26434 645289
rect 24899 644994 24905 645288
rect 25199 645284 26434 645288
rect 25199 644998 26143 645284
rect 26429 644998 26434 645284
rect 25199 644994 26434 644998
rect 24904 644993 26434 644994
rect 26778 645151 26948 645157
rect 26778 644993 26784 645151
rect 26942 644993 26948 645151
rect 26778 644987 26948 644993
rect 26365 644823 26687 644824
rect 26360 644503 26366 644823
rect 26686 644503 26692 644823
rect 26365 644502 26687 644503
rect 49828 643594 49834 643631
rect 7129 643298 24904 643594
rect 25200 643298 49834 643594
rect 50265 643594 50271 643631
rect 50265 643298 54241 643594
rect 7129 643202 7251 643298
rect 7469 643202 8723 643298
rect 8941 643202 10195 643298
rect 10413 643202 11667 643298
rect 11885 643202 13139 643298
rect 13357 643202 14611 643298
rect 14829 643202 16083 643298
rect 16301 643202 17555 643298
rect 17773 643202 19027 643298
rect 19245 643202 20499 643298
rect 20717 643202 21971 643298
rect 22189 643202 23443 643298
rect 23661 643202 24915 643298
rect 25133 643202 26387 643298
rect 26605 643202 27859 643298
rect 28077 643202 29331 643298
rect 29549 643202 30803 643298
rect 31021 643202 32275 643298
rect 32493 643202 33747 643298
rect 33965 643202 35219 643298
rect 35437 643202 36691 643298
rect 36909 643202 38163 643298
rect 38381 643202 39635 643298
rect 39853 643202 41107 643298
rect 41325 643202 42579 643298
rect 42797 643202 44051 643298
rect 44269 643202 45523 643298
rect 45741 643202 46995 643298
rect 47213 643202 48467 643298
rect 48685 643202 49834 643298
rect 50265 643202 51411 643298
rect 51629 643202 52883 643298
rect 53101 643202 54241 643298
rect 7129 643200 49834 643202
rect 50265 643200 54241 643202
rect 7129 643161 54241 643200
rect 7231 642755 54254 642763
rect 7231 642754 50444 642755
rect 7231 642658 7251 642754
rect 7469 642658 8723 642754
rect 8941 642658 10195 642754
rect 10413 642658 11667 642754
rect 11885 642658 13139 642754
rect 13357 642658 14611 642754
rect 14829 642658 16083 642754
rect 16301 642658 17555 642754
rect 17773 642658 19027 642754
rect 19245 642658 20499 642754
rect 20717 642658 21971 642754
rect 22189 642658 23443 642754
rect 23661 642658 24915 642754
rect 25133 642658 26387 642754
rect 26605 642658 27859 642754
rect 28077 642658 29331 642754
rect 29549 642658 30803 642754
rect 31021 642658 32275 642754
rect 32493 642658 33747 642754
rect 33965 642658 35219 642754
rect 35437 642658 36691 642754
rect 36909 642658 38163 642754
rect 38381 642658 39635 642754
rect 39853 642658 41107 642754
rect 41325 642658 42579 642754
rect 42797 642658 44051 642754
rect 44269 642658 45523 642754
rect 45741 642658 46995 642754
rect 47213 642658 48467 642754
rect 48685 642658 49939 642754
rect 50157 642658 50444 642754
rect 7231 642618 26365 642658
rect 7243 642336 26365 642618
rect 26687 642336 50444 642658
rect 50438 642330 50444 642336
rect 50869 642754 54254 642755
rect 50869 642658 51411 642754
rect 51629 642658 52883 642754
rect 53101 642658 54254 642754
rect 50869 642336 54254 642658
rect 50869 642330 50875 642336
rect 56264 641802 59030 642374
rect 56264 641577 57514 641802
rect 57739 641577 59030 641802
rect 5974 641447 8474 641551
rect 5974 641240 6999 641447
rect 7206 641240 8474 641447
rect -800 633842 1660 638642
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 5974 513753 8474 641240
rect 96 511642 8474 513753
rect -800 511530 8474 511642
rect 96 511253 8474 511530
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 5974 504876 8474 511253
rect 56264 470680 59030 641577
rect 582340 639784 584800 644584
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 245 468420 59030 470680
rect -800 468308 59030 468420
rect 245 467914 59030 468308
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect 126727 3535 127430 3540
rect 126726 3534 127431 3535
rect -800 2726 480 2838
rect 126726 2831 126727 3534
rect 127430 2831 127431 3534
rect 126726 2830 127431 2831
rect 126727 2825 127430 2830
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 173299 696988 175797 699486
rect 222483 699661 224981 702159
rect 324294 699894 326494 702094
rect 217176 696988 219674 699486
rect 413837 699895 416035 702093
rect 172231 691258 174731 693758
rect 49833 655930 50266 656363
rect 50443 653776 50870 654203
rect 24905 644994 25199 645288
rect 26784 645146 26942 645151
rect 26784 644998 26789 645146
rect 26789 644998 26937 645146
rect 26937 644998 26942 645146
rect 26784 644993 26942 644998
rect 26366 644819 26686 644823
rect 26366 644507 26370 644819
rect 26370 644507 26682 644819
rect 26682 644507 26686 644819
rect 26366 644503 26686 644507
rect 24904 643298 25200 643594
rect 49834 643298 50265 643631
rect 49834 643202 49939 643298
rect 49939 643202 50157 643298
rect 50157 643202 50265 643298
rect 49834 643200 50265 643202
rect 26365 642336 26687 642658
rect 50444 642330 50869 642755
rect 126727 3530 127430 3534
rect 126727 2835 126731 3530
rect 126731 2835 127426 3530
rect 127426 2835 127430 3530
rect 126727 2831 127430 2835
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702458 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 222482 702159 224982 702160
rect 222482 699661 222483 702159
rect 224981 699661 224982 702159
rect 324293 702094 326495 702095
rect 324293 699894 324294 702094
rect 326494 702093 416036 702094
rect 326494 699895 413837 702093
rect 416035 699895 416036 702093
rect 326494 699894 416036 699895
rect 324293 699893 326495 699894
rect 38828 699486 219675 699487
rect 38828 696988 173299 699486
rect 175797 696988 217176 699486
rect 219674 696988 219675 699486
rect 38828 696987 219675 696988
rect 38828 682040 41328 696987
rect 172230 693758 174732 693759
rect 222482 693758 224982 699661
rect 50678 691258 172231 693758
rect 174731 691258 224982 693758
rect 50678 679904 53178 691258
rect 172230 691257 174732 691258
rect 45260 677404 53178 679904
rect 49832 656363 50267 656364
rect 49832 655930 49833 656363
rect 50266 655930 50267 656363
rect 49832 655929 50267 655930
rect 24904 645288 25200 645289
rect 24904 644994 24905 645288
rect 25199 644994 25200 645288
rect 24904 643595 25200 644994
rect 26783 645151 26943 645152
rect 26783 644993 26784 645151
rect 26942 644993 26943 645151
rect 26783 644992 26943 644993
rect 26365 644823 26687 644824
rect 26365 644503 26366 644823
rect 26686 644503 26687 644823
rect 24903 643594 25201 643595
rect 24903 643298 24904 643594
rect 25200 643298 25201 643594
rect 24903 643297 25201 643298
rect 26365 642659 26687 644503
rect 26364 642658 26688 642659
rect 26364 642336 26365 642658
rect 26687 642336 26688 642658
rect 26364 642335 26688 642336
rect 26789 642084 26937 644992
rect 49833 643631 50266 655929
rect 50442 654203 50871 654204
rect 50442 653776 50443 654203
rect 50870 653776 50871 654203
rect 50442 653775 50871 653776
rect 49833 643200 49834 643631
rect 50265 643200 50266 643631
rect 49833 643199 50266 643200
rect 50443 642755 50870 653775
rect 50443 642330 50444 642755
rect 50869 642330 50870 642755
rect 50443 642329 50870 642330
rect 26789 642076 27418 642084
rect 26713 3535 27418 642076
rect 26713 3534 127431 3535
rect 26713 2831 126727 3534
rect 127430 2831 127431 3534
rect 26713 2830 127431 2831
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use cfg_shift_register  cfg_shift_register_0
timestamp 1646794523
transform 1 0 42470 0 1 642694
box -72 -183 11802 839
use cfg_shift_register  cfg_shift_register_1
timestamp 1646794523
transform 1 0 30694 0 1 642694
box -72 -183 11802 839
use cfg_shift_register  cfg_shift_register_2
timestamp 1646794523
transform 1 0 18918 0 1 642694
box -72 -183 11802 839
use cfg_shift_register  cfg_shift_register_3
timestamp 1646794523
transform 1 0 7142 0 1 642694
box -72 -183 11802 839
use proj_sstl_test  proj_sstl_test_0
timestamp 1646793240
transform 1 0 15929 0 1 645492
box -424 16 33306 40167
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646787781
transform 1 0 54234 0 1 642706
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1646787781
transform 1 0 7038 0 1 642706
box -38 -48 130 592
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
