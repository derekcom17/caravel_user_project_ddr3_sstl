magic
tech sky130A
magscale 1 2
timestamp 1646794523
<< nwell >>
rect -50 518 118 839
rect 5819 594 6350 646
rect 9819 594 10350 646
<< pwell >>
rect -9 -183 77 -26
<< psubdiff >>
rect 5905 -39 5939 -5
rect 5997 -39 6031 -5
rect 9905 -39 9939 -5
rect 9997 -39 10031 -5
rect 17 -99 51 -52
rect 17 -157 51 -133
<< nsubdiff >>
rect 17 771 51 795
rect 17 678 51 737
rect 17 620 51 644
rect 5905 573 5939 607
rect 5997 573 6031 607
rect 9905 573 9939 607
rect 9997 573 10031 607
<< psubdiffcont >>
rect 5939 -39 5997 -5
rect 9939 -39 9997 -5
rect 17 -133 51 -99
<< nsubdiffcont >>
rect 17 737 51 771
rect 17 644 51 678
rect 5939 573 5997 607
rect 9939 573 9997 607
<< locali >>
rect 5 771 63 806
rect 5 737 17 771
rect 51 737 63 771
rect 5 678 63 737
rect 5 644 17 678
rect 51 644 63 678
rect 5 573 63 644
rect 5923 573 5939 607
rect 5997 573 6013 607
rect 9923 573 9939 607
rect 9997 573 10013 607
rect -12 539 17 573
rect 51 539 80 573
rect -12 -5 17 29
rect 51 -5 80 29
rect 5 -99 63 -5
rect 5923 -39 5939 -5
rect 5997 -39 6013 -5
rect 9923 -39 9939 -5
rect 9997 -39 10013 -5
rect 5 -133 17 -99
rect 51 -133 63 -99
rect 5 -150 63 -133
<< viali >>
rect 17 539 51 573
rect 19 228 53 262
rect 1491 228 1525 262
rect 2963 228 2997 262
rect 4435 228 4469 262
rect 5907 228 5941 262
rect 7379 228 7413 262
rect 8851 228 8885 262
rect 10323 228 10357 262
rect 273 155 307 189
rect 1745 155 1779 189
rect 3217 155 3251 189
rect 4689 155 4723 189
rect 6161 155 6195 189
rect 7633 155 7667 189
rect 9105 155 9139 189
rect 10577 155 10611 189
rect 1370 101 1411 142
rect 2842 101 2883 142
rect 4314 101 4355 142
rect 5786 101 5827 142
rect 7258 101 7299 142
rect 8730 101 8771 142
rect 10202 101 10243 142
rect 11674 101 11715 142
rect 17 -5 51 29
<< metal1 >>
rect -12 573 80 604
rect -12 539 17 573
rect 51 539 80 573
rect -12 508 80 539
rect 7 267 65 268
rect 1479 267 1537 268
rect 2951 267 3009 268
rect 4423 267 4481 268
rect 5895 267 5953 268
rect 7367 267 7425 268
rect 8839 267 8897 268
rect 10311 267 10369 268
rect -60 262 11802 267
rect -60 228 19 262
rect 53 228 1491 262
rect 1525 228 2963 262
rect 2997 228 4435 262
rect 4469 228 5907 262
rect 5941 228 7379 262
rect 7413 228 8851 262
rect 8885 228 10323 262
rect 10357 228 11802 262
rect -60 223 11802 228
rect 7 222 65 223
rect 1479 222 1537 223
rect 2951 222 3009 223
rect 4423 222 4481 223
rect 5895 222 5953 223
rect 7367 222 7425 223
rect 8839 222 8897 223
rect 10311 222 10369 223
rect 236 189 319 195
rect 236 155 273 189
rect 307 155 319 189
rect -72 148 -14 154
rect -72 96 -66 148
rect 236 149 319 155
rect 1708 189 1791 195
rect 1708 155 1745 189
rect 1779 155 1791 189
rect 236 142 277 149
rect -14 101 277 142
rect 1364 148 1458 154
rect 1364 142 1406 148
rect 1708 149 1791 155
rect 3180 189 3263 195
rect 3180 155 3217 189
rect 3251 155 3263 189
rect 1708 142 1749 149
rect 1364 101 1370 142
rect 1458 101 1749 142
rect 2836 148 2930 154
rect 2836 142 2878 148
rect 3180 149 3263 155
rect 4652 189 4735 195
rect 4652 155 4689 189
rect 4723 155 4735 189
rect 3180 142 3221 149
rect 2836 101 2842 142
rect 2930 101 3221 142
rect 4308 148 4402 154
rect 4308 142 4350 148
rect 4652 149 4735 155
rect 6124 189 6207 195
rect 6124 155 6161 189
rect 6195 155 6207 189
rect 4652 142 4693 149
rect 4308 101 4314 142
rect 4402 101 4693 142
rect 5780 148 5874 154
rect 5780 142 5822 148
rect 6124 149 6207 155
rect 7596 189 7679 195
rect 7596 155 7633 189
rect 7667 155 7679 189
rect 6124 142 6165 149
rect 5780 101 5786 142
rect 5874 101 6165 142
rect 7252 148 7346 154
rect 7252 142 7294 148
rect 7596 149 7679 155
rect 9068 189 9151 195
rect 9068 155 9105 189
rect 9139 155 9151 189
rect 7596 142 7637 149
rect 7252 101 7258 142
rect 7346 101 7637 142
rect 8724 148 8818 154
rect 8724 142 8766 148
rect 9068 149 9151 155
rect 10540 189 10623 195
rect 10540 155 10577 189
rect 10611 155 10623 189
rect 9068 142 9109 149
rect 8724 101 8730 142
rect 8818 101 9109 142
rect 10196 148 10290 154
rect 10196 142 10238 148
rect 10540 149 10623 155
rect 10540 142 10581 149
rect 10196 101 10202 142
rect 10290 101 10581 142
rect 11668 148 11762 154
rect 11668 142 11710 148
rect 11668 101 11674 142
rect 11762 101 11802 142
rect -72 89 -14 96
rect 1364 96 1406 101
rect 1364 90 1458 96
rect 2836 96 2878 101
rect 2836 90 2930 96
rect 4308 96 4350 101
rect 4308 90 4402 96
rect 5780 96 5822 101
rect 5780 90 5874 96
rect 7252 96 7294 101
rect 7252 90 7346 96
rect 8724 96 8766 101
rect 8724 90 8818 96
rect 10196 96 10238 101
rect 10196 90 10290 96
rect 11668 96 11710 101
rect 11668 90 11762 96
rect 1364 89 1417 90
rect 2836 89 2889 90
rect 4308 89 4361 90
rect 5780 89 5833 90
rect 7252 89 7305 90
rect 8724 89 8777 90
rect 10196 89 10249 90
rect 11668 89 11721 90
rect -12 29 80 60
rect -12 -5 17 29
rect 51 -5 80 29
rect -12 -36 80 -5
<< via1 >>
rect -66 96 -14 148
rect 1406 142 1458 148
rect 1406 101 1411 142
rect 1411 101 1458 142
rect 2878 142 2930 148
rect 2878 101 2883 142
rect 2883 101 2930 142
rect 4350 142 4402 148
rect 4350 101 4355 142
rect 4355 101 4402 142
rect 5822 142 5874 148
rect 5822 101 5827 142
rect 5827 101 5874 142
rect 7294 142 7346 148
rect 7294 101 7299 142
rect 7299 101 7346 142
rect 8766 142 8818 148
rect 8766 101 8771 142
rect 8771 101 8818 142
rect 10238 142 10290 148
rect 10238 101 10243 142
rect 10243 101 10290 142
rect 11710 142 11762 148
rect 11710 101 11715 142
rect 11715 101 11762 142
rect 1406 96 1458 101
rect 2878 96 2930 101
rect 4350 96 4402 101
rect 5822 96 5874 101
rect 7294 96 7346 101
rect 8766 96 8818 101
rect 10238 96 10290 101
rect 11710 96 11762 101
<< metal2 >>
rect -60 148 -20 604
rect 1412 148 1452 604
rect 2884 148 2924 604
rect 4356 148 4396 604
rect 5828 148 5868 604
rect 7300 148 7340 604
rect 8772 148 8812 604
rect 10244 148 10284 604
rect 11716 148 11756 604
rect -72 96 -66 148
rect -14 96 -8 148
rect 1400 96 1406 148
rect 1458 96 1464 148
rect 2872 96 2878 148
rect 2930 96 2936 148
rect 4344 96 4350 148
rect 4402 96 4408 148
rect 5816 96 5822 148
rect 5874 96 5880 148
rect 7288 96 7294 148
rect 7346 96 7352 148
rect 8760 96 8766 148
rect 8818 96 8824 148
rect 10232 96 10238 148
rect 10290 96 10296 148
rect 11704 96 11710 148
rect 11762 96 11768 148
rect -60 -36 -20 96
rect 1412 -36 1452 96
rect 2884 -36 2924 96
rect 4356 -36 4396 96
rect 5828 -36 5868 96
rect 7300 -36 7340 96
rect 8772 -36 8812 96
rect 10244 -36 10284 96
rect 11716 -36 11756 96
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646794523
transform 1 0 -12 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1646794523
transform 1 0 1460 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1646794523
transform 1 0 2932 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1646794523
transform 1 0 4404 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1646794523
transform 1 0 5876 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1646794523
transform 1 0 7348 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1646794523
transform 1 0 8820 0 1 12
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1646794523
transform 1 0 10292 0 1 12
box -38 -48 1510 592
<< labels >>
flabel metal2 s -60 -36 -20 604 1 FreeSerif 480 0 0 0 d_in
port 1 n
flabel metal2 s 1412 -36 1452 604 1 FreeSerif 480 0 0 0 q[0]
port 3 n
flabel metal2 s 2884 -36 2924 604 1 FreeSerif 480 0 0 0 q[1]
port 4 n
flabel metal2 s 4356 -36 4396 604 1 FreeSerif 480 180 0 0 q[2]
port 5 n
flabel metal2 s 5828 -36 5868 604 1 FreeSerif 480 180 0 0 q[3]
port 6 n
flabel metal2 s 7300 -36 7340 604 1 FreeSerif 480 180 0 0 q[4]
port 7 n
flabel metal2 s 8772 -36 8812 604 1 FreeSerif 480 180 0 0 q[5]
port 8 n
flabel metal2 s 10244 -36 10284 604 1 FreeSerif 480 180 0 0 q[6]
port 9 n
flabel metal2 s 11716 -36 11756 604 1 FreeSerif 480 180 0 0 q[7]
port 10 n
flabel metal1 s 10357 223 11802 267 1 FreeSerif 480 0 0 0 clk
port 0 n
flabel metal1 s -12 508 80 604 1 FreeSerif 320 0 0 0 VDD
port 11 n
flabel metal1 s -12 -36 80 60 1 FreeSerif 320 0 0 0 GND
port 2 n
<< end >>
