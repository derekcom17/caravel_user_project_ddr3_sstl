* NGSPICE file created from SSTL.ext - technology: sky130A

.subckt n-leg_ctrl_fet_2 a_n125_n65# a_n81_n153# a_n33_n65# VSUBS
X0 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=4.03e+11p ps=3.84e+06u w=650000u l=150000u
X1 a_n33_n65# a_n81_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n125_n65# a_n81_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt n-leg_ctrl_fet_0 a_n125_n153# a_n125_n65# a_n33_n65# VSUBS
X0 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=3.4255e+12p pd=3.264e+07u as=3.432e+12p ps=3.136e+07u w=650000u l=150000u
X1 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt n-leg_ctrl_fet_3 a_15_n19# a_n73_n19# a_n33_n107# VSUBS
X0 a_15_n19# a_n33_n107# a_n73_n19# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt n-leg_ctrl_fet_1 a_n125_n153# a_n125_n65# a_n33_n65# VSUBS
X0 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=7.84e+06u as=1.0075e+12p ps=9.6e+06u w=650000u l=150000u
X1 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_n33_n65# a_n125_n153# a_n125_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_n125_n65# a_n125_n153# a_n33_n65# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt n-leg_polyres a_n33_170# a_n33_n243#
R0 a_n33_n243# a_n33_170# sky130_fd_pr__res_generic_po w=330000u l=1.7e+06u
.ends

.subckt n-leg pd_ctrl DQ cal_ctrl[0] cal_ctrl[1] cal_ctrl[2] cal_ctrl[3] li_1854_527#
+ GND
Xn-leg_ctrl_fet_2_0 DQ cal_ctrl[2] vpulldown GND n-leg_ctrl_fet_2
Xn-leg_ctrl_fet_0_0 cal_ctrl[0] DQ vpulldown GND n-leg_ctrl_fet_0
Xn-leg_ctrl_fet_3_0 DQ vpulldown cal_ctrl[3] GND n-leg_ctrl_fet_3
Xn-leg_ctrl_fet_1_0 cal_ctrl[1] vpulldown DQ GND n-leg_ctrl_fet_1
Xn-leg_polyres_0 vpulldown DQ n-leg_polyres
X0 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=1.20215e+13p pd=2.595e+06u as=9.6163e+12p ps=9.0425e+07u w=650000u l=150000u
X1 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X42 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 GND pd_ctrl vpulldown GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt p-leg_fet_16 a_n1053_n161# a_n1053_n64# a_995_n64# a_n285_n64# a_n541_n64#
+ a_483_n64# a_739_n64# a_n29_n64# a_n925_n64# a_227_n64# w_n1089_n100# a_n797_n64#
X0 a_n925_n64# a_n1053_n161# a_n541_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n797_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X2 a_n925_n64# a_n1053_n161# a_227_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X3 a_739_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X4 a_n925_n64# a_n1053_n161# a_n29_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_n285_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X6 a_n925_n64# a_n1053_n161# a_n797_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X7 a_227_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X8 a_n925_n64# a_n1053_n161# a_483_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X9 a_995_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X10 a_n925_n64# a_n1053_n161# a_n1053_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X11 a_n925_n64# a_n1053_n161# a_739_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X12 a_n541_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X13 a_n925_n64# a_n1053_n161# a_n285_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X14 a_n29_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X15 a_483_n64# a_n1053_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt p-leg_polyres a_n33_n253# a_n33_180#
R0 a_n33_n253# a_n33_180# sky130_fd_pr__res_generic_po w=330000u l=1.8e+06u
.ends

.subckt p-leg_6 a_n1053_n64# a_n285_n64# a_n541_n64# a_n995_n161# a_n925_n64# w_n1089_n100#
+ a_n797_n64#
X0 a_n925_n64# a_n995_n161# a_n541_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n797_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X2 a_n285_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X3 a_n925_n64# a_n995_n161# a_n797_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X4 a_n925_n64# a_n995_n161# a_n1053_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_n541_n64# a_n995_n161# a_n925_n64# w_n1089_n100# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt p-leg DQ VDD n_cal_ctrl[0] n_cal_ctrl[1] n_cal_ctrl[2] n_cal_ctrl[3] n_pu_ctrl
+ w_3710_2162# li_4_2169# w_1502_2162# w_4446_2162# w_2974_2162# w_2238_2162# w_5918_2162#
+ extr_sky130_fd_sc_hd__fill_8_9/VPWR w_766_2162# extr_sky130_fd_sc_hd__fill_8_8/VGND extr_sky130_fd_sc_hd__fill_8_9/VGND
+ w_5182_2162#
Xp-leg_fet_16_4 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
Xp-leg_fet_16_5 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
Xp-leg_fet_16_6 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_fet_16
Xp-leg_fet_16_7 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_fet_16
Xp-leg_polyres_0 DQ li_16_1957# p-leg_polyres
Xp-leg_fet_16_8 n_cal_ctrl[0] li_16_1957# li_16_1957# li_16_1957# li_16_1957# li_16_1957#
+ li_16_1957# li_16_1957# DQ li_16_1957# VDD li_16_1957# p-leg_fet_16
Xp-leg_6_0 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6
Xp-leg_6_1 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6
Xp-leg_6_2 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6
Xp-leg_6_3 DQ DQ DQ n_cal_ctrl[1] li_16_1957# VDD DQ p-leg_6
Xp-leg_6_4 DQ DQ DQ n_cal_ctrl[2] li_16_1957# VDD DQ p-leg_6
Xp-leg_6_6 li_16_1957# li_16_1957# li_16_1957# n_cal_ctrl[3] DQ VDD li_16_1957# p-leg_6
Xp-leg_6_5 DQ DQ DQ n_cal_ctrl[2] li_16_1957# VDD DQ p-leg_6
Xp-leg_fet_16_0 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
Xp-leg_fet_16_1 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
Xp-leg_fet_16_2 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
Xp-leg_fet_16_3 n_pu_ctrl VDD VDD VDD VDD VDD VDD VDD li_16_1957# VDD VDD VDD p-leg_fet_16
.ends

.subckt extr_sky130_fd_sc_hd__clkbuf_8 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=6.951e+11p ps=8.35e+06u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt extr_sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt extr_sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt extr_sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt extr_sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt SSTL DQ GND pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3] pd_ctrl[0]
+ pd_ctrl[1] pd_ctrl[2] pd_ctrl[3] pd_ctrl[4] pd_ctrl[5] pd_ctrl[6] pu_cal_ctrl[0]
+ pu_cal_ctrl[1] pu_cal_ctrl[2] pu_cal_ctrl[3] pu_ctrl[0] pu_ctrl[1] pu_ctrl[2] pu_ctrl[3]
+ pu_ctrl[4] pu_ctrl[5] pu_ctrl[6] VDD
Xn-leg_0 n-leg_0/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xp-leg_3 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_3/n_pu_ctrl p-leg_3/w_3710_2162# GND p-leg_3/w_1502_2162#
+ p-leg_3/w_4446_2162# p-leg_3/w_2974_2162# p-leg_3/w_2238_2162# p-leg_3/w_5918_2162#
+ p-leg_3/extr_sky130_fd_sc_hd__fill_8_9/VPWR p-leg_3/w_766_2162# GND GND p-leg_3/w_5182_2162#
+ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_1 extr_sky130_fd_sc_hd__clkinv_4_2/Y GND VDD n-leg_1/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xn-leg_1 n-leg_1/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xp-leg_4 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_4/n_pu_ctrl p-leg_4/w_3710_2162# GND p-leg_4/w_1502_2162#
+ p-leg_4/w_4446_2162# p-leg_4/w_2974_2162# p-leg_4/w_2238_2162# p-leg_4/w_5918_2162#
+ p-leg_4/extr_sky130_fd_sc_hd__fill_8_9/VPWR p-leg_4/w_766_2162# GND GND p-leg_4/w_5182_2162#
+ p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_2 extr_sky130_fd_sc_hd__clkinv_4_4/Y GND VDD n-leg_2/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xn-leg_2 n-leg_2/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xp-leg_5 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_5/n_pu_ctrl p-leg_5/w_3710_2162# GND p-leg_5/w_1502_2162#
+ p-leg_5/w_4446_2162# p-leg_5/w_2974_2162# p-leg_5/w_2238_2162# p-leg_5/w_5918_2162#
+ VDD p-leg_5/w_766_2162# GND GND p-leg_5/w_5182_2162# p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_3 extr_sky130_fd_sc_hd__clkinv_4_6/Y GND VDD n-leg_3/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_10 extr_sky130_fd_sc_hd__clkinv_4_11/Y GND VDD extr_sky130_fd_sc_hd__clkbuf_8_5/A
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_3 n-leg_3/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xp-leg_6 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_6/n_pu_ctrl p-leg_6/w_3710_2162# GND p-leg_6/w_1502_2162#
+ p-leg_6/w_4446_2162# p-leg_6/w_2974_2162# p-leg_6/w_2238_2162# p-leg_6/w_5918_2162#
+ p-leg_6/extr_sky130_fd_sc_hd__fill_8_9/VPWR p-leg_6/w_766_2162# GND GND p-leg_6/w_5182_2162#
+ p-leg
Xextr_sky130_fd_sc_hd__clkinv_16_0 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_4 extr_sky130_fd_sc_hd__clkinv_4_8/Y GND VDD n-leg_4/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_11 pd_ctrl[5] GND VDD extr_sky130_fd_sc_hd__clkinv_4_11/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_4 n-leg_4/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_16_1 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_5 extr_sky130_fd_sc_hd__clkbuf_8_5/A GND VDD n-leg_5/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_12 extr_sky130_fd_sc_hd__clkinv_4_13/Y GND VDD extr_sky130_fd_sc_hd__clkbuf_8_6/A
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_5 n-leg_5/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_16_2 extr_sky130_fd_sc_hd__clkinv_16_2/A GND VDD p-leg_0/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_8_6 extr_sky130_fd_sc_hd__clkbuf_8_6/A GND VDD n-leg_6/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
Xextr_sky130_fd_sc_hd__clkinv_4_13 pd_ctrl[6] GND VDD extr_sky130_fd_sc_hd__clkinv_4_13/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xn-leg_6 n-leg_6/pd_ctrl DQ pd_cal_ctrl[0] pd_cal_ctrl[1] pd_cal_ctrl[2] pd_cal_ctrl[3]
+ VDD GND n-leg
Xextr_sky130_fd_sc_hd__clkinv_4_0 extr_sky130_fd_sc_hd__clkinv_4_1/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_0/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_3 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_1 pd_ctrl[0] GND VDD extr_sky130_fd_sc_hd__clkinv_4_1/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_4 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_2 extr_sky130_fd_sc_hd__clkinv_4_3/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_2/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_5 extr_sky130_fd_sc_hd__clkinv_16_5/A GND VDD p-leg_1/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_3 pd_ctrl[1] GND VDD extr_sky130_fd_sc_hd__clkinv_4_3/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_6 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_4 extr_sky130_fd_sc_hd__clkinv_4_5/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_4/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_7 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_5 pd_ctrl[2] GND VDD extr_sky130_fd_sc_hd__clkinv_4_5/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_8 extr_sky130_fd_sc_hd__clkinv_16_8/A GND VDD p-leg_2/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_20 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_6 extr_sky130_fd_sc_hd__clkinv_4_7/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_6/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_9 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_10 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_7 pd_ctrl[3] GND VDD extr_sky130_fd_sc_hd__clkinv_4_7/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_4_8 extr_sky130_fd_sc_hd__clkinv_4_9/Y GND VDD extr_sky130_fd_sc_hd__clkinv_4_8/Y
+ GND VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_11 extr_sky130_fd_sc_hd__clkinv_16_9/A GND VDD p-leg_3/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_12 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_4_9 pd_ctrl[4] GND VDD extr_sky130_fd_sc_hd__clkinv_4_9/Y GND
+ VDD extr_sky130_fd_sc_hd__clkinv_4
Xextr_sky130_fd_sc_hd__clkinv_16_13 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_14 extr_sky130_fd_sc_hd__clkbuf_16_4/X GND VDD p-leg_4/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_15 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkinv_16_16 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_0 pu_ctrl[0] GND VDD extr_sky130_fd_sc_hd__clkinv_16_2/A GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_17 extr_sky130_fd_sc_hd__clkbuf_16_5/X GND VDD p-leg_5/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_1 pu_ctrl[1] GND VDD extr_sky130_fd_sc_hd__clkinv_16_5/A GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_18 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_2 pu_ctrl[2] GND VDD extr_sky130_fd_sc_hd__clkinv_16_8/A GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkinv_16_19 extr_sky130_fd_sc_hd__clkbuf_16_6/X GND VDD p-leg_6/n_pu_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkinv_16
Xextr_sky130_fd_sc_hd__clkbuf_16_3 pu_ctrl[3] GND VDD extr_sky130_fd_sc_hd__clkinv_16_9/A GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_4 pu_ctrl[4] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_4/X GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_5 pu_ctrl[5] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_5/X GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__clkbuf_16_6 pu_ctrl[6] GND VDD extr_sky130_fd_sc_hd__clkbuf_16_6/X GND
+ VDD extr_sky130_fd_sc_hd__clkbuf_16
Xextr_sky130_fd_sc_hd__inv_1_0 pu_cal_ctrl[0] GND VDD p-leg_6/n_cal_ctrl[0] GND VDD extr_sky130_fd_sc_hd__inv_1
Xextr_sky130_fd_sc_hd__inv_1_1 pu_cal_ctrl[1] GND VDD p-leg_6/n_cal_ctrl[1] GND VDD extr_sky130_fd_sc_hd__inv_1
Xp-leg_0 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_0/n_pu_ctrl GND GND GND GND GND GND GND p-leg_0/extr_sky130_fd_sc_hd__fill_8_9/VPWR
+ GND GND GND GND p-leg
Xp-leg_1 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_1/n_pu_ctrl p-leg_1/w_3710_2162# GND p-leg_1/w_1502_2162#
+ p-leg_1/w_4446_2162# p-leg_1/w_2974_2162# p-leg_1/w_2238_2162# p-leg_1/w_5918_2162#
+ p-leg_1/extr_sky130_fd_sc_hd__fill_8_9/VPWR p-leg_1/w_766_2162# GND GND p-leg_1/w_5182_2162#
+ p-leg
Xextr_sky130_fd_sc_hd__inv_1_2 pu_cal_ctrl[2] GND VDD p-leg_6/n_cal_ctrl[2] GND VDD extr_sky130_fd_sc_hd__inv_1
Xextr_sky130_fd_sc_hd__inv_1_3 pu_cal_ctrl[3] GND VDD p-leg_6/n_cal_ctrl[3] GND VDD extr_sky130_fd_sc_hd__inv_1
Xp-leg_2 DQ VDD p-leg_6/n_cal_ctrl[0] p-leg_6/n_cal_ctrl[1] p-leg_6/n_cal_ctrl[2]
+ p-leg_6/n_cal_ctrl[3] p-leg_2/n_pu_ctrl p-leg_2/w_3710_2162# GND p-leg_2/w_1502_2162#
+ p-leg_2/w_4446_2162# p-leg_2/w_2974_2162# p-leg_2/w_2238_2162# p-leg_2/w_5918_2162#
+ VDD p-leg_2/w_766_2162# GND GND p-leg_2/w_5182_2162# p-leg
Xextr_sky130_fd_sc_hd__clkbuf_8_0 extr_sky130_fd_sc_hd__clkinv_4_0/Y GND VDD n-leg_0/pd_ctrl
+ GND VDD extr_sky130_fd_sc_hd__clkbuf_8
.ends

