// SPDX-FileCopyrightText: 2020 University of Washingington CSE
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
`timescale 1 ns / 1 ps

/*
   TODO add description
*/

module cfg_shift_register (
    input clk,    // Clock
    input din, // Clock Enable
    output [0:31] q
);

    always @(posedge clk) begin
        q[1:31] <= q[0:30];
        q[0] <= din;
    end

endmodule