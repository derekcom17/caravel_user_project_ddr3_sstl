magic
tech sky130A
magscale 1 2
timestamp 1646874728
<< error_p >>
rect -125 -65 -63 65
rect -33 -65 33 65
rect 63 -65 125 65
rect 155 -65 221 65
<< nmos >>
rect -63 -65 -33 65
rect 33 -65 63 65
rect 125 -65 155 65
<< ndiff >>
rect -125 57 -63 65
rect -125 17 -113 57
rect -79 17 -63 57
rect -125 -65 -63 17
rect -33 -17 33 65
rect -33 -57 -17 -17
rect 17 -57 33 -17
rect -33 -65 33 -57
rect 63 57 125 65
rect 63 17 75 57
rect 109 17 125 57
rect 63 -65 125 17
rect 155 -17 221 65
rect 155 -57 171 -17
rect 205 -57 221 -17
rect 155 -65 221 -57
<< ndiffc >>
rect -113 17 -79 57
rect -17 -57 17 -17
rect 75 17 109 57
rect 171 -57 205 -17
<< poly >>
rect -63 65 -33 91
rect 33 65 63 91
rect 125 65 155 91
rect -63 -87 -33 -65
rect 33 -87 63 -65
rect 125 -87 155 -65
rect -81 -103 173 -87
rect -81 -137 -65 -103
rect -31 -137 31 -103
rect 65 -137 123 -103
rect 157 -137 173 -103
rect -81 -153 173 -137
<< polycont >>
rect -65 -137 -31 -103
rect 31 -137 65 -103
rect 123 -137 157 -103
<< locali >>
rect -129 17 -113 57
rect -79 17 75 57
rect 109 17 221 57
rect -129 -57 -17 -17
rect 17 -57 171 -17
rect 205 -57 221 -17
rect -81 -137 -65 -103
rect -31 -137 31 -103
rect 65 -137 123 -103
rect 157 -137 173 -103
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.650 l 0.150 m 1 nf 2 diffcov 25 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
