magic
tech sky130A
magscale 1 2
timestamp 1646875043
<< pwell >>
rect 1883 1071 1917 1105
rect 3355 1071 3389 1105
rect 4827 1071 4861 1105
rect 1854 21 3314 203
rect 3340 21 4786 203
rect 4812 21 6258 203
rect 1883 -17 1917 21
rect 3355 -17 3389 21
rect 4827 -17 4861 21
<< scnmos >>
rect 1946 47 1976 177
rect 2030 47 2060 177
rect 2114 47 2144 177
rect 2198 47 2228 177
rect 2282 47 2312 177
rect 2366 47 2396 177
rect 2450 47 2480 177
rect 2534 47 2564 177
rect 2618 47 2648 177
rect 2702 47 2732 177
rect 2786 47 2816 177
rect 2870 47 2900 177
rect 2954 47 2984 177
rect 3038 47 3068 177
rect 3122 47 3152 177
rect 3206 47 3236 177
rect 3418 47 3448 177
rect 3502 47 3532 177
rect 3586 47 3616 177
rect 3670 47 3700 177
rect 3754 47 3784 177
rect 3838 47 3868 177
rect 3922 47 3952 177
rect 4006 47 4036 177
rect 4090 47 4120 177
rect 4174 47 4204 177
rect 4258 47 4288 177
rect 4342 47 4372 177
rect 4426 47 4456 177
rect 4510 47 4540 177
rect 4594 47 4624 177
rect 4678 47 4708 177
rect 4890 47 4920 177
rect 4974 47 5004 177
rect 5058 47 5088 177
rect 5142 47 5172 177
rect 5226 47 5256 177
rect 5310 47 5340 177
rect 5394 47 5424 177
rect 5478 47 5508 177
rect 5562 47 5592 177
rect 5646 47 5676 177
rect 5730 47 5760 177
rect 5814 47 5844 177
rect 5898 47 5928 177
rect 5982 47 6012 177
rect 6066 47 6096 177
rect 6150 47 6180 177
<< ndiff >>
rect 6325 808 6361 812
rect 6325 782 6331 808
rect 1864 161 1946 177
rect 1864 127 1902 161
rect 1936 127 1946 161
rect 1864 93 1946 127
rect 1864 59 1902 93
rect 1936 59 1946 93
rect 1864 47 1946 59
rect 1976 161 2030 177
rect 1976 127 1986 161
rect 2020 127 2030 161
rect 1976 93 2030 127
rect 1976 59 1986 93
rect 2020 59 2030 93
rect 1976 47 2030 59
rect 2060 93 2114 177
rect 2060 59 2070 93
rect 2104 59 2114 93
rect 2060 47 2114 59
rect 2144 161 2198 177
rect 2144 127 2154 161
rect 2188 127 2198 161
rect 2144 93 2198 127
rect 2144 59 2154 93
rect 2188 59 2198 93
rect 2144 47 2198 59
rect 2228 93 2282 177
rect 2228 59 2238 93
rect 2272 59 2282 93
rect 2228 47 2282 59
rect 2312 161 2366 177
rect 2312 127 2322 161
rect 2356 127 2366 161
rect 2312 93 2366 127
rect 2312 59 2322 93
rect 2356 59 2366 93
rect 2312 47 2366 59
rect 2396 93 2450 177
rect 2396 59 2406 93
rect 2440 59 2450 93
rect 2396 47 2450 59
rect 2480 161 2534 177
rect 2480 127 2490 161
rect 2524 127 2534 161
rect 2480 93 2534 127
rect 2480 59 2490 93
rect 2524 59 2534 93
rect 2480 47 2534 59
rect 2564 93 2618 177
rect 2564 59 2574 93
rect 2608 59 2618 93
rect 2564 47 2618 59
rect 2648 161 2702 177
rect 2648 127 2658 161
rect 2692 127 2702 161
rect 2648 93 2702 127
rect 2648 59 2658 93
rect 2692 59 2702 93
rect 2648 47 2702 59
rect 2732 93 2786 177
rect 2732 59 2742 93
rect 2776 59 2786 93
rect 2732 47 2786 59
rect 2816 161 2870 177
rect 2816 127 2826 161
rect 2860 127 2870 161
rect 2816 93 2870 127
rect 2816 59 2826 93
rect 2860 59 2870 93
rect 2816 47 2870 59
rect 2900 93 2954 177
rect 2900 59 2910 93
rect 2944 59 2954 93
rect 2900 47 2954 59
rect 2984 161 3038 177
rect 2984 127 2994 161
rect 3028 127 3038 161
rect 2984 93 3038 127
rect 2984 59 2994 93
rect 3028 59 3038 93
rect 2984 47 3038 59
rect 3068 93 3122 177
rect 3068 59 3078 93
rect 3112 59 3122 93
rect 3068 47 3122 59
rect 3152 161 3206 177
rect 3152 127 3162 161
rect 3196 127 3206 161
rect 3152 93 3206 127
rect 3152 59 3162 93
rect 3196 59 3206 93
rect 3152 47 3206 59
rect 3236 161 3288 177
rect 3236 127 3246 161
rect 3280 127 3288 161
rect 3236 93 3288 127
rect 3236 59 3246 93
rect 3280 59 3288 93
rect 3236 47 3288 59
rect 3366 161 3418 177
rect 3366 127 3374 161
rect 3408 127 3418 161
rect 3366 93 3418 127
rect 3366 59 3374 93
rect 3408 59 3418 93
rect 3366 47 3418 59
rect 3448 161 3502 177
rect 3448 127 3458 161
rect 3492 127 3502 161
rect 3448 93 3502 127
rect 3448 59 3458 93
rect 3492 59 3502 93
rect 3448 47 3502 59
rect 3532 93 3586 177
rect 3532 59 3542 93
rect 3576 59 3586 93
rect 3532 47 3586 59
rect 3616 161 3670 177
rect 3616 127 3626 161
rect 3660 127 3670 161
rect 3616 93 3670 127
rect 3616 59 3626 93
rect 3660 59 3670 93
rect 3616 47 3670 59
rect 3700 93 3754 177
rect 3700 59 3710 93
rect 3744 59 3754 93
rect 3700 47 3754 59
rect 3784 161 3838 177
rect 3784 127 3794 161
rect 3828 127 3838 161
rect 3784 93 3838 127
rect 3784 59 3794 93
rect 3828 59 3838 93
rect 3784 47 3838 59
rect 3868 93 3922 177
rect 3868 59 3878 93
rect 3912 59 3922 93
rect 3868 47 3922 59
rect 3952 161 4006 177
rect 3952 127 3962 161
rect 3996 127 4006 161
rect 3952 93 4006 127
rect 3952 59 3962 93
rect 3996 59 4006 93
rect 3952 47 4006 59
rect 4036 93 4090 177
rect 4036 59 4046 93
rect 4080 59 4090 93
rect 4036 47 4090 59
rect 4120 161 4174 177
rect 4120 127 4130 161
rect 4164 127 4174 161
rect 4120 93 4174 127
rect 4120 59 4130 93
rect 4164 59 4174 93
rect 4120 47 4174 59
rect 4204 93 4258 177
rect 4204 59 4214 93
rect 4248 59 4258 93
rect 4204 47 4258 59
rect 4288 161 4342 177
rect 4288 127 4298 161
rect 4332 127 4342 161
rect 4288 93 4342 127
rect 4288 59 4298 93
rect 4332 59 4342 93
rect 4288 47 4342 59
rect 4372 93 4426 177
rect 4372 59 4382 93
rect 4416 59 4426 93
rect 4372 47 4426 59
rect 4456 161 4510 177
rect 4456 127 4466 161
rect 4500 127 4510 161
rect 4456 93 4510 127
rect 4456 59 4466 93
rect 4500 59 4510 93
rect 4456 47 4510 59
rect 4540 93 4594 177
rect 4540 59 4550 93
rect 4584 59 4594 93
rect 4540 47 4594 59
rect 4624 161 4678 177
rect 4624 127 4634 161
rect 4668 127 4678 161
rect 4624 93 4678 127
rect 4624 59 4634 93
rect 4668 59 4678 93
rect 4624 47 4678 59
rect 4708 161 4760 177
rect 4708 127 4718 161
rect 4752 127 4760 161
rect 4708 93 4760 127
rect 4708 59 4718 93
rect 4752 59 4760 93
rect 4708 47 4760 59
rect 4838 161 4890 177
rect 4838 127 4846 161
rect 4880 127 4890 161
rect 4838 93 4890 127
rect 4838 59 4846 93
rect 4880 59 4890 93
rect 4838 47 4890 59
rect 4920 161 4974 177
rect 4920 127 4930 161
rect 4964 127 4974 161
rect 4920 93 4974 127
rect 4920 59 4930 93
rect 4964 59 4974 93
rect 4920 47 4974 59
rect 5004 93 5058 177
rect 5004 59 5014 93
rect 5048 59 5058 93
rect 5004 47 5058 59
rect 5088 161 5142 177
rect 5088 127 5098 161
rect 5132 127 5142 161
rect 5088 93 5142 127
rect 5088 59 5098 93
rect 5132 59 5142 93
rect 5088 47 5142 59
rect 5172 93 5226 177
rect 5172 59 5182 93
rect 5216 59 5226 93
rect 5172 47 5226 59
rect 5256 161 5310 177
rect 5256 127 5266 161
rect 5300 127 5310 161
rect 5256 93 5310 127
rect 5256 59 5266 93
rect 5300 59 5310 93
rect 5256 47 5310 59
rect 5340 93 5394 177
rect 5340 59 5350 93
rect 5384 59 5394 93
rect 5340 47 5394 59
rect 5424 161 5478 177
rect 5424 127 5434 161
rect 5468 127 5478 161
rect 5424 93 5478 127
rect 5424 59 5434 93
rect 5468 59 5478 93
rect 5424 47 5478 59
rect 5508 93 5562 177
rect 5508 59 5518 93
rect 5552 59 5562 93
rect 5508 47 5562 59
rect 5592 161 5646 177
rect 5592 127 5602 161
rect 5636 127 5646 161
rect 5592 93 5646 127
rect 5592 59 5602 93
rect 5636 59 5646 93
rect 5592 47 5646 59
rect 5676 93 5730 177
rect 5676 59 5686 93
rect 5720 59 5730 93
rect 5676 47 5730 59
rect 5760 161 5814 177
rect 5760 127 5770 161
rect 5804 127 5814 161
rect 5760 93 5814 127
rect 5760 59 5770 93
rect 5804 59 5814 93
rect 5760 47 5814 59
rect 5844 93 5898 177
rect 5844 59 5854 93
rect 5888 59 5898 93
rect 5844 47 5898 59
rect 5928 161 5982 177
rect 5928 127 5938 161
rect 5972 127 5982 161
rect 5928 93 5982 127
rect 5928 59 5938 93
rect 5972 59 5982 93
rect 5928 47 5982 59
rect 6012 93 6066 177
rect 6012 59 6022 93
rect 6056 59 6066 93
rect 6012 47 6066 59
rect 6096 161 6150 177
rect 6096 127 6106 161
rect 6140 127 6150 161
rect 6096 93 6150 127
rect 6096 59 6106 93
rect 6140 59 6150 93
rect 6096 47 6150 59
rect 6180 161 6232 177
rect 6180 127 6190 161
rect 6224 127 6232 161
rect 6180 93 6232 127
rect 6180 59 6190 93
rect 6224 59 6232 93
rect 6180 47 6232 59
<< ndiffc >>
rect 1902 127 1936 161
rect 1902 59 1936 93
rect 1986 127 2020 161
rect 1986 59 2020 93
rect 2070 59 2104 93
rect 2154 127 2188 161
rect 2154 59 2188 93
rect 2238 59 2272 93
rect 2322 127 2356 161
rect 2322 59 2356 93
rect 2406 59 2440 93
rect 2490 127 2524 161
rect 2490 59 2524 93
rect 2574 59 2608 93
rect 2658 127 2692 161
rect 2658 59 2692 93
rect 2742 59 2776 93
rect 2826 127 2860 161
rect 2826 59 2860 93
rect 2910 59 2944 93
rect 2994 127 3028 161
rect 2994 59 3028 93
rect 3078 59 3112 93
rect 3162 127 3196 161
rect 3162 59 3196 93
rect 3246 127 3280 161
rect 3246 59 3280 93
rect 3374 127 3408 161
rect 3374 59 3408 93
rect 3458 127 3492 161
rect 3458 59 3492 93
rect 3542 59 3576 93
rect 3626 127 3660 161
rect 3626 59 3660 93
rect 3710 59 3744 93
rect 3794 127 3828 161
rect 3794 59 3828 93
rect 3878 59 3912 93
rect 3962 127 3996 161
rect 3962 59 3996 93
rect 4046 59 4080 93
rect 4130 127 4164 161
rect 4130 59 4164 93
rect 4214 59 4248 93
rect 4298 127 4332 161
rect 4298 59 4332 93
rect 4382 59 4416 93
rect 4466 127 4500 161
rect 4466 59 4500 93
rect 4550 59 4584 93
rect 4634 127 4668 161
rect 4634 59 4668 93
rect 4718 127 4752 161
rect 4718 59 4752 93
rect 4846 127 4880 161
rect 4846 59 4880 93
rect 4930 127 4964 161
rect 4930 59 4964 93
rect 5014 59 5048 93
rect 5098 127 5132 161
rect 5098 59 5132 93
rect 5182 59 5216 93
rect 5266 127 5300 161
rect 5266 59 5300 93
rect 5350 59 5384 93
rect 5434 127 5468 161
rect 5434 59 5468 93
rect 5518 59 5552 93
rect 5602 127 5636 161
rect 5602 59 5636 93
rect 5686 59 5720 93
rect 5770 127 5804 161
rect 5770 59 5804 93
rect 5854 59 5888 93
rect 5938 127 5972 161
rect 5938 59 5972 93
rect 6022 59 6056 93
rect 6106 127 6140 161
rect 6106 59 6140 93
rect 6190 127 6224 161
rect 6190 59 6224 93
<< psubdiff >>
rect 1975 1071 2009 1105
rect 2067 1071 2101 1105
rect 6286 156 6519 180
rect 6286 21 6519 45
<< psubdiffcont >>
rect 2009 1071 2067 1105
rect 6286 45 6519 156
<< poly >>
rect 1854 249 6270 265
rect 1854 215 1950 249
rect 1984 215 2070 249
rect 2104 215 2238 249
rect 2272 215 2407 249
rect 2441 215 2574 249
rect 2608 215 2742 249
rect 2776 215 2909 249
rect 2943 215 3076 249
rect 3110 215 3243 249
rect 3277 215 3368 249
rect 3402 215 3542 249
rect 3576 215 3710 249
rect 3744 215 3879 249
rect 3913 215 4046 249
rect 4080 215 4214 249
rect 4248 215 4381 249
rect 4415 215 4548 249
rect 4582 215 4715 249
rect 4749 215 4840 249
rect 4874 215 5014 249
rect 5048 215 5182 249
rect 5216 215 5351 249
rect 5385 215 5518 249
rect 5552 215 5686 249
rect 5720 215 5853 249
rect 5887 215 6020 249
rect 6054 215 6187 249
rect 6221 215 6270 249
rect 1854 199 6270 215
rect 1946 177 1976 199
rect 2030 177 2060 199
rect 2114 177 2144 199
rect 2198 177 2228 199
rect 2282 177 2312 199
rect 2366 177 2396 199
rect 2450 177 2480 199
rect 2534 177 2564 199
rect 2618 177 2648 199
rect 2702 177 2732 199
rect 2786 177 2816 199
rect 2870 177 2900 199
rect 2954 177 2984 199
rect 3038 177 3068 199
rect 3122 177 3152 199
rect 3206 177 3236 199
rect 3418 177 3448 199
rect 3502 177 3532 199
rect 3586 177 3616 199
rect 3670 177 3700 199
rect 3754 177 3784 199
rect 3838 177 3868 199
rect 3922 177 3952 199
rect 4006 177 4036 199
rect 4090 177 4120 199
rect 4174 177 4204 199
rect 4258 177 4288 199
rect 4342 177 4372 199
rect 4426 177 4456 199
rect 4510 177 4540 199
rect 4594 177 4624 199
rect 4678 177 4708 199
rect 4890 177 4920 199
rect 4974 177 5004 199
rect 5058 177 5088 199
rect 5142 177 5172 199
rect 5226 177 5256 199
rect 5310 177 5340 199
rect 5394 177 5424 199
rect 5478 177 5508 199
rect 5562 177 5592 199
rect 5646 177 5676 199
rect 5730 177 5760 199
rect 5814 177 5844 199
rect 5898 177 5928 199
rect 5982 177 6012 199
rect 6066 177 6096 199
rect 6150 177 6180 199
rect 1946 21 1976 47
rect 2030 21 2060 47
rect 2114 21 2144 47
rect 2198 21 2228 47
rect 2282 21 2312 47
rect 2366 21 2396 47
rect 2450 21 2480 47
rect 2534 21 2564 47
rect 2618 21 2648 47
rect 2702 21 2732 47
rect 2786 21 2816 47
rect 2870 21 2900 47
rect 2954 21 2984 47
rect 3038 21 3068 47
rect 3122 21 3152 47
rect 3206 21 3236 47
rect 3418 21 3448 47
rect 3502 21 3532 47
rect 3586 21 3616 47
rect 3670 21 3700 47
rect 3754 21 3784 47
rect 3838 21 3868 47
rect 3922 21 3952 47
rect 4006 21 4036 47
rect 4090 21 4120 47
rect 4174 21 4204 47
rect 4258 21 4288 47
rect 4342 21 4372 47
rect 4426 21 4456 47
rect 4510 21 4540 47
rect 4594 21 4624 47
rect 4678 21 4708 47
rect 4890 21 4920 47
rect 4974 21 5004 47
rect 5058 21 5088 47
rect 5142 21 5172 47
rect 5226 21 5256 47
rect 5310 21 5340 47
rect 5394 21 5424 47
rect 5478 21 5508 47
rect 5562 21 5592 47
rect 5646 21 5676 47
rect 5730 21 5760 47
rect 5814 21 5844 47
rect 5898 21 5928 47
rect 5982 21 6012 47
rect 6066 21 6096 47
rect 6150 21 6180 47
<< polycont >>
rect 1950 215 1984 249
rect 2070 215 2104 249
rect 2238 215 2272 249
rect 2407 215 2441 249
rect 2574 215 2608 249
rect 2742 215 2776 249
rect 2909 215 2943 249
rect 3076 215 3110 249
rect 3243 215 3277 249
rect 3368 215 3402 249
rect 3542 215 3576 249
rect 3710 215 3744 249
rect 3879 215 3913 249
rect 4046 215 4080 249
rect 4214 215 4248 249
rect 4381 215 4415 249
rect 4548 215 4582 249
rect 4715 215 4749 249
rect 4840 215 4874 249
rect 5014 215 5048 249
rect 5182 215 5216 249
rect 5351 215 5385 249
rect 5518 215 5552 249
rect 5686 215 5720 249
rect 5853 215 5887 249
rect 6020 215 6054 249
rect 6187 215 6221 249
<< locali >>
rect 1854 1071 1883 1105
rect 1917 1071 1975 1105
rect 2101 1071 2159 1105
rect 2193 1071 2251 1105
rect 2285 1071 2343 1105
rect 2377 1071 2435 1105
rect 2469 1071 2527 1105
rect 2561 1071 2619 1105
rect 2653 1071 2711 1105
rect 2745 1071 2803 1105
rect 2837 1071 2895 1105
rect 2929 1071 2987 1105
rect 3021 1071 3079 1105
rect 3113 1071 3171 1105
rect 3205 1071 3263 1105
rect 3297 1071 3355 1105
rect 3389 1071 3447 1105
rect 3481 1071 3539 1105
rect 3573 1071 3631 1105
rect 3665 1071 3723 1105
rect 3757 1071 3815 1105
rect 3849 1071 3907 1105
rect 3941 1071 3999 1105
rect 4033 1071 4091 1105
rect 4125 1071 4183 1105
rect 4217 1071 4275 1105
rect 4309 1071 4367 1105
rect 4401 1071 4459 1105
rect 4493 1071 4551 1105
rect 4585 1071 4643 1105
rect 4677 1071 4735 1105
rect 4769 1071 4827 1105
rect 4861 1071 4919 1105
rect 4953 1071 5011 1105
rect 5045 1071 5103 1105
rect 5137 1071 5195 1105
rect 5229 1071 5287 1105
rect 5321 1071 5379 1105
rect 5413 1071 5471 1105
rect 5505 1071 5563 1105
rect 5597 1071 5655 1105
rect 5689 1071 5747 1105
rect 5781 1071 5839 1105
rect 5873 1071 5931 1105
rect 5965 1071 6023 1105
rect 6057 1071 6115 1105
rect 6149 1071 6207 1105
rect 6241 1071 6299 1105
rect 6333 1071 6391 1105
rect 6425 1071 6483 1105
rect 6517 1071 6546 1105
rect 4936 886 5004 926
rect 4970 852 5004 886
rect 5887 864 6023 904
rect 6325 864 6465 904
rect 5887 852 5921 864
rect 4970 812 5039 852
rect 5853 812 5921 852
rect 4902 778 4936 812
rect 5955 790 6019 830
rect 6325 812 6377 830
rect 6431 812 6465 864
rect 6325 790 6363 812
rect 5955 778 5989 790
rect 4902 738 5039 778
rect 5853 738 5989 778
rect 1854 527 1883 561
rect 1917 527 1975 561
rect 2009 527 2067 561
rect 2101 527 2159 561
rect 2193 527 2251 561
rect 2285 527 2343 561
rect 2377 527 2435 561
rect 2469 527 2527 561
rect 2561 527 2619 561
rect 2653 527 2711 561
rect 2745 527 2803 561
rect 2837 527 2895 561
rect 2929 527 2987 561
rect 3021 527 3079 561
rect 3113 527 3171 561
rect 3205 527 3263 561
rect 3297 527 3355 561
rect 3389 527 3447 561
rect 3481 527 3539 561
rect 3573 527 3631 561
rect 3665 527 3723 561
rect 3757 527 3815 561
rect 3849 527 3907 561
rect 3941 527 3999 561
rect 4033 527 4091 561
rect 4125 527 4183 561
rect 4217 527 4275 561
rect 4309 527 4367 561
rect 4401 527 4459 561
rect 4493 527 4551 561
rect 4585 527 4643 561
rect 4677 527 4735 561
rect 4769 527 4827 561
rect 4861 527 4919 561
rect 4953 527 5011 561
rect 5045 527 5103 561
rect 5137 527 5195 561
rect 5229 527 5287 561
rect 5321 527 5379 561
rect 5413 527 5471 561
rect 5505 527 5563 561
rect 5597 527 5655 561
rect 5689 527 5747 561
rect 5781 527 5839 561
rect 5873 527 5931 561
rect 5965 527 6023 561
rect 6057 527 6115 561
rect 6149 527 6207 561
rect 6241 527 6299 561
rect 6333 527 6391 561
rect 6425 527 6483 561
rect 6517 527 6546 561
rect 1854 249 6270 263
rect 1854 215 1950 249
rect 1984 215 2070 249
rect 2104 215 2238 249
rect 2272 215 2407 249
rect 2441 215 2574 249
rect 2608 215 2742 249
rect 2776 215 2909 249
rect 2943 215 3076 249
rect 3110 215 3243 249
rect 3277 215 3368 249
rect 3402 215 3542 249
rect 3576 215 3710 249
rect 3744 215 3879 249
rect 3913 215 4046 249
rect 4080 215 4214 249
rect 4248 215 4381 249
rect 4415 215 4548 249
rect 4582 215 4715 249
rect 4749 215 4840 249
rect 4874 215 5014 249
rect 5048 215 5182 249
rect 5216 215 5351 249
rect 5385 215 5518 249
rect 5552 215 5686 249
rect 5720 215 5853 249
rect 5887 215 6020 249
rect 6054 215 6187 249
rect 6221 215 6270 249
rect 1970 179 3212 181
rect 1890 161 1936 177
rect 1890 127 1902 161
rect 1890 93 1936 127
rect 1890 59 1902 93
rect 1890 17 1936 59
rect 1970 161 2069 179
rect 1970 127 1986 161
rect 2020 145 2069 161
rect 2103 161 2237 179
rect 2103 145 2154 161
rect 2020 143 2154 145
rect 2020 127 2036 143
rect 1970 93 2036 127
rect 2138 127 2154 143
rect 2188 145 2237 161
rect 2271 161 2405 179
rect 2271 145 2322 161
rect 2188 143 2322 145
rect 2188 127 2204 143
rect 1970 59 1986 93
rect 2020 59 2036 93
rect 1970 51 2036 59
rect 2070 93 2104 109
rect 2070 17 2104 59
rect 2138 93 2204 127
rect 2306 127 2322 143
rect 2356 145 2405 161
rect 2439 161 2573 179
rect 2439 145 2490 161
rect 2356 143 2490 145
rect 2356 127 2372 143
rect 2138 59 2154 93
rect 2188 59 2204 93
rect 2138 51 2204 59
rect 2238 93 2272 109
rect 2238 17 2272 59
rect 2306 93 2372 127
rect 2474 127 2490 143
rect 2524 145 2573 161
rect 2607 161 2741 179
rect 2607 145 2658 161
rect 2524 143 2658 145
rect 2524 127 2540 143
rect 2306 59 2322 93
rect 2356 59 2372 93
rect 2306 51 2372 59
rect 2406 93 2440 109
rect 2406 17 2440 59
rect 2474 93 2540 127
rect 2642 127 2658 143
rect 2692 145 2741 161
rect 2775 161 2909 179
rect 2775 145 2826 161
rect 2692 143 2826 145
rect 2692 127 2708 143
rect 2474 59 2490 93
rect 2524 59 2540 93
rect 2474 51 2540 59
rect 2574 93 2608 109
rect 2574 17 2608 59
rect 2642 93 2708 127
rect 2810 127 2826 143
rect 2860 145 2909 161
rect 2943 161 3077 179
rect 2943 145 2994 161
rect 2860 143 2994 145
rect 2860 127 2876 143
rect 2642 59 2658 93
rect 2692 59 2708 93
rect 2642 51 2708 59
rect 2742 93 2776 109
rect 2742 17 2776 59
rect 2810 93 2876 127
rect 2978 127 2994 143
rect 3028 145 3077 161
rect 3111 161 3212 179
rect 3442 179 4684 181
rect 3111 145 3162 161
rect 3028 143 3162 145
rect 3028 127 3044 143
rect 2810 59 2826 93
rect 2860 59 2876 93
rect 2810 51 2876 59
rect 2910 93 2944 109
rect 2910 17 2944 59
rect 2978 93 3044 127
rect 3146 127 3162 143
rect 3196 127 3212 161
rect 2978 59 2994 93
rect 3028 59 3044 93
rect 2978 51 3044 59
rect 3078 93 3112 109
rect 3078 17 3112 59
rect 3146 93 3212 127
rect 3146 59 3162 93
rect 3196 59 3212 93
rect 3146 51 3212 59
rect 3246 161 3288 177
rect 3280 127 3288 161
rect 3246 93 3288 127
rect 3280 59 3288 93
rect 3246 17 3288 59
rect 3362 161 3408 177
rect 3362 127 3374 161
rect 3362 93 3408 127
rect 3362 59 3374 93
rect 3362 17 3408 59
rect 3442 161 3541 179
rect 3442 127 3458 161
rect 3492 145 3541 161
rect 3575 161 3709 179
rect 3575 145 3626 161
rect 3492 143 3626 145
rect 3492 127 3508 143
rect 3442 93 3508 127
rect 3610 127 3626 143
rect 3660 145 3709 161
rect 3743 161 3877 179
rect 3743 145 3794 161
rect 3660 143 3794 145
rect 3660 127 3676 143
rect 3442 59 3458 93
rect 3492 59 3508 93
rect 3442 51 3508 59
rect 3542 93 3576 109
rect 3542 17 3576 59
rect 3610 93 3676 127
rect 3778 127 3794 143
rect 3828 145 3877 161
rect 3911 161 4045 179
rect 3911 145 3962 161
rect 3828 143 3962 145
rect 3828 127 3844 143
rect 3610 59 3626 93
rect 3660 59 3676 93
rect 3610 51 3676 59
rect 3710 93 3744 109
rect 3710 17 3744 59
rect 3778 93 3844 127
rect 3946 127 3962 143
rect 3996 145 4045 161
rect 4079 161 4213 179
rect 4079 145 4130 161
rect 3996 143 4130 145
rect 3996 127 4012 143
rect 3778 59 3794 93
rect 3828 59 3844 93
rect 3778 51 3844 59
rect 3878 93 3912 109
rect 3878 17 3912 59
rect 3946 93 4012 127
rect 4114 127 4130 143
rect 4164 145 4213 161
rect 4247 161 4381 179
rect 4247 145 4298 161
rect 4164 143 4298 145
rect 4164 127 4180 143
rect 3946 59 3962 93
rect 3996 59 4012 93
rect 3946 51 4012 59
rect 4046 93 4080 109
rect 4046 17 4080 59
rect 4114 93 4180 127
rect 4282 127 4298 143
rect 4332 145 4381 161
rect 4415 161 4549 179
rect 4415 145 4466 161
rect 4332 143 4466 145
rect 4332 127 4348 143
rect 4114 59 4130 93
rect 4164 59 4180 93
rect 4114 51 4180 59
rect 4214 93 4248 109
rect 4214 17 4248 59
rect 4282 93 4348 127
rect 4450 127 4466 143
rect 4500 145 4549 161
rect 4583 161 4684 179
rect 4914 179 6156 181
rect 4583 145 4634 161
rect 4500 143 4634 145
rect 4500 127 4516 143
rect 4282 59 4298 93
rect 4332 59 4348 93
rect 4282 51 4348 59
rect 4382 93 4416 109
rect 4382 17 4416 59
rect 4450 93 4516 127
rect 4618 127 4634 143
rect 4668 127 4684 161
rect 4450 59 4466 93
rect 4500 59 4516 93
rect 4450 51 4516 59
rect 4550 93 4584 109
rect 4550 17 4584 59
rect 4618 93 4684 127
rect 4618 59 4634 93
rect 4668 59 4684 93
rect 4618 51 4684 59
rect 4718 161 4760 177
rect 4752 127 4760 161
rect 4718 93 4760 127
rect 4752 59 4760 93
rect 4718 17 4760 59
rect 4834 161 4880 177
rect 4834 127 4846 161
rect 4834 93 4880 127
rect 4834 59 4846 93
rect 4834 17 4880 59
rect 4914 161 5013 179
rect 4914 127 4930 161
rect 4964 145 5013 161
rect 5047 161 5181 179
rect 5047 145 5098 161
rect 4964 143 5098 145
rect 4964 127 4980 143
rect 4914 93 4980 127
rect 5082 127 5098 143
rect 5132 145 5181 161
rect 5215 161 5349 179
rect 5215 145 5266 161
rect 5132 143 5266 145
rect 5132 127 5148 143
rect 4914 59 4930 93
rect 4964 59 4980 93
rect 4914 51 4980 59
rect 5014 93 5048 109
rect 5014 17 5048 59
rect 5082 93 5148 127
rect 5250 127 5266 143
rect 5300 145 5349 161
rect 5383 161 5517 179
rect 5383 145 5434 161
rect 5300 143 5434 145
rect 5300 127 5316 143
rect 5082 59 5098 93
rect 5132 59 5148 93
rect 5082 51 5148 59
rect 5182 93 5216 109
rect 5182 17 5216 59
rect 5250 93 5316 127
rect 5418 127 5434 143
rect 5468 145 5517 161
rect 5551 161 5685 179
rect 5551 145 5602 161
rect 5468 143 5602 145
rect 5468 127 5484 143
rect 5250 59 5266 93
rect 5300 59 5316 93
rect 5250 51 5316 59
rect 5350 93 5384 109
rect 5350 17 5384 59
rect 5418 93 5484 127
rect 5586 127 5602 143
rect 5636 145 5685 161
rect 5719 161 5853 179
rect 5719 145 5770 161
rect 5636 143 5770 145
rect 5636 127 5652 143
rect 5418 59 5434 93
rect 5468 59 5484 93
rect 5418 51 5484 59
rect 5518 93 5552 109
rect 5518 17 5552 59
rect 5586 93 5652 127
rect 5754 127 5770 143
rect 5804 145 5853 161
rect 5887 161 6021 179
rect 5887 145 5938 161
rect 5804 143 5938 145
rect 5804 127 5820 143
rect 5586 59 5602 93
rect 5636 59 5652 93
rect 5586 51 5652 59
rect 5686 93 5720 109
rect 5686 17 5720 59
rect 5754 93 5820 127
rect 5922 127 5938 143
rect 5972 145 6021 161
rect 6055 161 6156 179
rect 6055 145 6106 161
rect 5972 143 6106 145
rect 5972 127 5988 143
rect 5754 59 5770 93
rect 5804 59 5820 93
rect 5754 51 5820 59
rect 5854 93 5888 109
rect 5854 17 5888 59
rect 5922 93 5988 127
rect 6090 127 6106 143
rect 6140 127 6156 161
rect 5922 59 5938 93
rect 5972 59 5988 93
rect 5922 51 5988 59
rect 6022 93 6056 109
rect 6022 17 6056 59
rect 6090 93 6156 127
rect 6090 59 6106 93
rect 6140 59 6156 93
rect 6090 51 6156 59
rect 6190 161 6232 177
rect 6224 127 6232 161
rect 6190 93 6232 127
rect 6224 59 6232 93
rect 6190 17 6232 59
rect 6286 156 6519 180
rect 6286 17 6519 45
rect 1854 -17 1883 17
rect 1917 -17 1975 17
rect 2009 -17 2067 17
rect 2101 -17 2159 17
rect 2193 -17 2251 17
rect 2285 -17 2343 17
rect 2377 -17 2435 17
rect 2469 -17 2527 17
rect 2561 -17 2619 17
rect 2653 -17 2711 17
rect 2745 -17 2803 17
rect 2837 -17 2895 17
rect 2929 -17 2987 17
rect 3021 -17 3079 17
rect 3113 -17 3171 17
rect 3205 -17 3263 17
rect 3297 -17 3355 17
rect 3389 -17 3447 17
rect 3481 -17 3539 17
rect 3573 -17 3631 17
rect 3665 -17 3723 17
rect 3757 -17 3815 17
rect 3849 -17 3907 17
rect 3941 -17 3999 17
rect 4033 -17 4091 17
rect 4125 -17 4183 17
rect 4217 -17 4275 17
rect 4309 -17 4367 17
rect 4401 -17 4459 17
rect 4493 -17 4551 17
rect 4585 -17 4643 17
rect 4677 -17 4735 17
rect 4769 -17 4827 17
rect 4861 -17 4919 17
rect 4953 -17 5011 17
rect 5045 -17 5103 17
rect 5137 -17 5195 17
rect 5229 -17 5287 17
rect 5321 -17 5379 17
rect 5413 -17 5471 17
rect 5505 -17 5563 17
rect 5597 -17 5655 17
rect 5689 -17 5747 17
rect 5781 -17 5839 17
rect 5873 -17 5931 17
rect 5965 -17 6023 17
rect 6057 -17 6115 17
rect 6149 -17 6207 17
rect 6241 -17 6299 17
rect 6333 -17 6391 17
rect 6425 -17 6483 17
rect 6517 -17 6546 17
<< viali >>
rect 1883 1071 1917 1105
rect 1975 1071 2009 1105
rect 2067 1071 2101 1105
rect 2159 1071 2193 1105
rect 2251 1071 2285 1105
rect 2343 1071 2377 1105
rect 2435 1071 2469 1105
rect 2527 1071 2561 1105
rect 2619 1071 2653 1105
rect 2711 1071 2745 1105
rect 2803 1071 2837 1105
rect 2895 1071 2929 1105
rect 2987 1071 3021 1105
rect 3079 1071 3113 1105
rect 3171 1071 3205 1105
rect 3263 1071 3297 1105
rect 3355 1071 3389 1105
rect 3447 1071 3481 1105
rect 3539 1071 3573 1105
rect 3631 1071 3665 1105
rect 3723 1071 3757 1105
rect 3815 1071 3849 1105
rect 3907 1071 3941 1105
rect 3999 1071 4033 1105
rect 4091 1071 4125 1105
rect 4183 1071 4217 1105
rect 4275 1071 4309 1105
rect 4367 1071 4401 1105
rect 4459 1071 4493 1105
rect 4551 1071 4585 1105
rect 4643 1071 4677 1105
rect 4735 1071 4769 1105
rect 4827 1071 4861 1105
rect 4919 1071 4953 1105
rect 5011 1071 5045 1105
rect 5103 1071 5137 1105
rect 5195 1071 5229 1105
rect 5287 1071 5321 1105
rect 5379 1071 5413 1105
rect 5471 1071 5505 1105
rect 5563 1071 5597 1105
rect 5655 1071 5689 1105
rect 5747 1071 5781 1105
rect 5839 1071 5873 1105
rect 5931 1071 5965 1105
rect 6023 1071 6057 1105
rect 6115 1071 6149 1105
rect 6207 1071 6241 1105
rect 6299 1071 6333 1105
rect 6391 1071 6425 1105
rect 6483 1071 6517 1105
rect 1866 972 4880 1006
rect 3980 886 4076 926
rect 5039 898 5853 932
rect 4426 812 4522 852
rect 6023 710 6277 744
rect 6371 636 6437 670
rect 1883 527 1917 561
rect 1975 527 2009 561
rect 2067 527 2101 561
rect 2159 527 2193 561
rect 2251 527 2285 561
rect 2343 527 2377 561
rect 2435 527 2469 561
rect 2527 527 2561 561
rect 2619 527 2653 561
rect 2711 527 2745 561
rect 2803 527 2837 561
rect 2895 527 2929 561
rect 2987 527 3021 561
rect 3079 527 3113 561
rect 3171 527 3205 561
rect 3263 527 3297 561
rect 3355 527 3389 561
rect 3447 527 3481 561
rect 3539 527 3573 561
rect 3631 527 3665 561
rect 3723 527 3757 561
rect 3815 527 3849 561
rect 3907 527 3941 561
rect 3999 527 4033 561
rect 4091 527 4125 561
rect 4183 527 4217 561
rect 4275 527 4309 561
rect 4367 527 4401 561
rect 4459 527 4493 561
rect 4551 527 4585 561
rect 4643 527 4677 561
rect 4735 527 4769 561
rect 4827 527 4861 561
rect 4919 527 4953 561
rect 5011 527 5045 561
rect 5103 527 5137 561
rect 5195 527 5229 561
rect 5287 527 5321 561
rect 5379 527 5413 561
rect 5471 527 5505 561
rect 5563 527 5597 561
rect 5655 527 5689 561
rect 5747 527 5781 561
rect 5839 527 5873 561
rect 5931 527 5965 561
rect 6023 527 6057 561
rect 6115 527 6149 561
rect 6207 527 6241 561
rect 6299 527 6333 561
rect 6391 527 6425 561
rect 6483 527 6517 561
rect 2069 145 2103 179
rect 2237 145 2271 179
rect 2405 145 2439 179
rect 2573 145 2607 179
rect 2741 145 2775 179
rect 2909 145 2943 179
rect 3077 145 3111 179
rect 3541 145 3575 179
rect 3709 145 3743 179
rect 3877 145 3911 179
rect 4045 145 4079 179
rect 4213 145 4247 179
rect 4381 145 4415 179
rect 4549 145 4583 179
rect 5013 145 5047 179
rect 5181 145 5215 179
rect 5349 145 5383 179
rect 5517 145 5551 179
rect 5685 145 5719 179
rect 5853 145 5887 179
rect 6021 145 6055 179
rect 1883 -17 1917 17
rect 1975 -17 2009 17
rect 2067 -17 2101 17
rect 2159 -17 2193 17
rect 2251 -17 2285 17
rect 2343 -17 2377 17
rect 2435 -17 2469 17
rect 2527 -17 2561 17
rect 2619 -17 2653 17
rect 2711 -17 2745 17
rect 2803 -17 2837 17
rect 2895 -17 2929 17
rect 2987 -17 3021 17
rect 3079 -17 3113 17
rect 3171 -17 3205 17
rect 3263 -17 3297 17
rect 3355 -17 3389 17
rect 3447 -17 3481 17
rect 3539 -17 3573 17
rect 3631 -17 3665 17
rect 3723 -17 3757 17
rect 3815 -17 3849 17
rect 3907 -17 3941 17
rect 3999 -17 4033 17
rect 4091 -17 4125 17
rect 4183 -17 4217 17
rect 4275 -17 4309 17
rect 4367 -17 4401 17
rect 4459 -17 4493 17
rect 4551 -17 4585 17
rect 4643 -17 4677 17
rect 4735 -17 4769 17
rect 4827 -17 4861 17
rect 4919 -17 4953 17
rect 5011 -17 5045 17
rect 5103 -17 5137 17
rect 5195 -17 5229 17
rect 5287 -17 5321 17
rect 5379 -17 5413 17
rect 5471 -17 5505 17
rect 5563 -17 5597 17
rect 5655 -17 5689 17
rect 5747 -17 5781 17
rect 5839 -17 5873 17
rect 5931 -17 5965 17
rect 6023 -17 6057 17
rect 6115 -17 6149 17
rect 6207 -17 6241 17
rect 6299 -17 6333 17
rect 6391 -17 6425 17
rect 6483 -17 6517 17
<< metal1 >>
rect 1854 1105 6546 1136
rect 1854 1071 1883 1105
rect 1917 1071 1975 1105
rect 2009 1071 2067 1105
rect 2101 1071 2159 1105
rect 2193 1071 2251 1105
rect 2285 1071 2343 1105
rect 2377 1071 2435 1105
rect 2469 1071 2527 1105
rect 2561 1071 2619 1105
rect 2653 1071 2711 1105
rect 2745 1071 2803 1105
rect 2837 1071 2895 1105
rect 2929 1071 2987 1105
rect 3021 1071 3079 1105
rect 3113 1071 3171 1105
rect 3205 1071 3263 1105
rect 3297 1071 3355 1105
rect 3389 1071 3447 1105
rect 3481 1071 3539 1105
rect 3573 1071 3631 1105
rect 3665 1071 3723 1105
rect 3757 1071 3815 1105
rect 3849 1071 3907 1105
rect 3941 1071 3999 1105
rect 4033 1071 4091 1105
rect 4125 1071 4183 1105
rect 4217 1071 4275 1105
rect 4309 1071 4367 1105
rect 4401 1071 4459 1105
rect 4493 1071 4551 1105
rect 4585 1071 4643 1105
rect 4677 1071 4735 1105
rect 4769 1071 4827 1105
rect 4861 1071 4919 1105
rect 4953 1071 5011 1105
rect 5045 1071 5103 1105
rect 5137 1071 5195 1105
rect 5229 1071 5287 1105
rect 5321 1071 5379 1105
rect 5413 1071 5471 1105
rect 5505 1071 5563 1105
rect 5597 1071 5655 1105
rect 5689 1071 5747 1105
rect 5781 1071 5839 1105
rect 5873 1071 5931 1105
rect 5965 1071 6023 1105
rect 6057 1071 6115 1105
rect 6149 1071 6207 1105
rect 6241 1071 6299 1105
rect 6333 1071 6391 1105
rect 6425 1071 6483 1105
rect 6517 1071 6546 1105
rect 1854 1040 6546 1071
rect 1854 1006 6546 1012
rect 1854 972 1866 1006
rect 4880 972 6546 1006
rect 1854 966 6546 972
rect 4227 932 5935 938
rect 3974 926 3980 932
rect 4076 926 4082 932
rect 1854 880 3566 926
rect 3968 886 3980 926
rect 4076 886 4088 926
rect 4227 898 5039 932
rect 5853 926 5935 932
rect 5853 898 6546 926
rect 4227 892 6546 898
rect 3974 880 3980 886
rect 4076 880 4082 886
rect 3520 824 3566 880
rect 4227 824 4273 892
rect 5889 880 6546 892
rect 4420 852 4426 858
rect 4522 852 4528 858
rect 3520 778 4273 824
rect 4414 812 4426 852
rect 4522 812 4534 852
rect 4420 806 4426 812
rect 4522 806 4528 812
rect 1854 744 6546 750
rect 1854 710 6023 744
rect 6277 710 6546 744
rect 1854 704 6546 710
rect 1854 670 6546 676
rect 1854 636 6371 670
rect 6437 636 6546 670
rect 1854 630 6546 636
rect 1854 561 6546 592
rect 1854 527 1883 561
rect 1917 527 1975 561
rect 2009 527 2067 561
rect 2101 527 2159 561
rect 2193 527 2251 561
rect 2285 527 2343 561
rect 2377 527 2435 561
rect 2469 527 2527 561
rect 2561 527 2619 561
rect 2653 527 2711 561
rect 2745 527 2803 561
rect 2837 527 2895 561
rect 2929 527 2987 561
rect 3021 527 3079 561
rect 3113 527 3171 561
rect 3205 527 3263 561
rect 3297 527 3355 561
rect 3389 527 3447 561
rect 3481 527 3539 561
rect 3573 527 3631 561
rect 3665 527 3723 561
rect 3757 527 3815 561
rect 3849 527 3907 561
rect 3941 527 3999 561
rect 4033 527 4091 561
rect 4125 527 4183 561
rect 4217 527 4275 561
rect 4309 527 4367 561
rect 4401 527 4459 561
rect 4493 527 4551 561
rect 4585 527 4643 561
rect 4677 527 4735 561
rect 4769 527 4827 561
rect 4861 527 4919 561
rect 4953 527 5011 561
rect 5045 527 5103 561
rect 5137 527 5195 561
rect 5229 527 5287 561
rect 5321 527 5379 561
rect 5413 527 5471 561
rect 5505 527 5563 561
rect 5597 527 5655 561
rect 5689 527 5747 561
rect 5781 527 5839 561
rect 5873 527 5931 561
rect 5965 527 6023 561
rect 6057 527 6115 561
rect 6149 527 6207 561
rect 6241 527 6299 561
rect 6333 527 6391 561
rect 6425 527 6483 561
rect 6517 527 6546 561
rect 1854 496 6546 527
rect 3980 431 4076 445
rect 3980 379 3999 431
rect 4051 379 4076 431
rect 3980 349 4076 379
rect 4426 412 4593 421
rect 4426 360 4438 412
rect 4490 360 4593 412
rect 4426 210 4593 360
rect 1854 179 6270 210
rect 1854 145 2069 179
rect 2103 145 2237 179
rect 2271 145 2405 179
rect 2439 145 2573 179
rect 2607 145 2741 179
rect 2775 145 2909 179
rect 2943 145 3077 179
rect 3111 145 3541 179
rect 3575 145 3709 179
rect 3743 145 3877 179
rect 3911 145 4045 179
rect 4079 145 4213 179
rect 4247 145 4381 179
rect 4415 145 4549 179
rect 4583 145 5013 179
rect 5047 145 5181 179
rect 5215 145 5349 179
rect 5383 145 5517 179
rect 5551 145 5685 179
rect 5719 145 5853 179
rect 5887 145 6021 179
rect 6055 145 6270 179
rect 1854 114 6270 145
rect 1854 17 6546 48
rect 1854 -17 1883 17
rect 1917 -17 1975 17
rect 2009 -17 2067 17
rect 2101 -17 2159 17
rect 2193 -17 2251 17
rect 2285 -17 2343 17
rect 2377 -17 2435 17
rect 2469 -17 2527 17
rect 2561 -17 2619 17
rect 2653 -17 2711 17
rect 2745 -17 2803 17
rect 2837 -17 2895 17
rect 2929 -17 2987 17
rect 3021 -17 3079 17
rect 3113 -17 3171 17
rect 3205 -17 3263 17
rect 3297 -17 3355 17
rect 3389 -17 3447 17
rect 3481 -17 3539 17
rect 3573 -17 3631 17
rect 3665 -17 3723 17
rect 3757 -17 3815 17
rect 3849 -17 3907 17
rect 3941 -17 3999 17
rect 4033 -17 4091 17
rect 4125 -17 4183 17
rect 4217 -17 4275 17
rect 4309 -17 4367 17
rect 4401 -17 4459 17
rect 4493 -17 4551 17
rect 4585 -17 4643 17
rect 4677 -17 4735 17
rect 4769 -17 4827 17
rect 4861 -17 4919 17
rect 4953 -17 5011 17
rect 5045 -17 5103 17
rect 5137 -17 5195 17
rect 5229 -17 5287 17
rect 5321 -17 5379 17
rect 5413 -17 5471 17
rect 5505 -17 5563 17
rect 5597 -17 5655 17
rect 5689 -17 5747 17
rect 5781 -17 5839 17
rect 5873 -17 5931 17
rect 5965 -17 6023 17
rect 6057 -17 6115 17
rect 6149 -17 6207 17
rect 6241 -17 6299 17
rect 6333 -17 6391 17
rect 6425 -17 6483 17
rect 6517 -17 6546 17
rect 1854 -48 6546 -17
<< via1 >>
rect 3980 926 4076 932
rect 3980 886 4076 926
rect 3980 880 4076 886
rect 4426 852 4522 858
rect 4426 812 4522 852
rect 4426 806 4522 812
rect 3999 379 4051 431
rect 4438 360 4490 412
<< metal2 >>
rect 3980 932 4076 938
rect 3980 431 4076 880
rect 3980 379 3999 431
rect 4051 379 4076 431
rect 3980 349 4076 379
rect 4426 858 4522 864
rect 4426 412 4522 806
rect 4426 360 4438 412
rect 4490 360 4522 412
rect 4426 349 4522 360
use n-leg_ctrl_fet_0  n-leg_ctrl_fet_0_0
timestamp 1646874728
transform 1 0 1991 0 -1 869
box -129 -153 2945 91
use n-leg_ctrl_fet_1  n-leg_ctrl_fet_1_0
timestamp 1646874728
transform 1 0 5164 0 -1 795
box -129 -153 689 91
use n-leg_ctrl_fet_2  n-leg_ctrl_fet_2_0
timestamp 1646874728
transform 1 0 6104 0 1 847
box -129 -153 221 91
use n-leg_ctrl_fet_3  n-leg_ctrl_fet_3_0
timestamp 1646874728
transform 1 0 6404 0 1 727
box -73 -107 73 107
use n-leg_polyres  n-leg_polyres_0
timestamp 1642386543
transform 0 1 4251 -1 0 398
box -33 -243 33 243
<< labels >>
flabel metal1 1900 733 1900 733 7 FreeSerif 320 0 0 0 cal_ctrl[2]
port 7 w
flabel metal1 1900 651 1900 651 7 FreeSerif 320 0 0 0 cal_ctrl[3]
port 8 w
flabel viali 1900 -1 1900 -1 7 FreeSerif 320 0 0 0 GND
port 2 w
flabel viali 1900 1089 1900 1089 7 FreeSerif 320 0 0 0 GND
port 2 w
flabel metal1 s 1900 995 1900 995 7 FreeSerif 320 0 0 0 cal_ctrl[0]
port 5 w
flabel metal2 4033 370 4033 370 7 FreeSerif 320 0 0 0 DQ
port 3 w
flabel metal1 s 1900 909 1900 909 7 FreeSerif 320 0 0 0 cal_ctrl[1]
port 6 w
flabel polycont 1967 232 1967 232 7 FreeSerif 320 0 0 0 pd_ctrl
port 1 w
<< end >>
