magic
tech sky130A
magscale 1 2
timestamp 1644116513
<< nwell >>
rect 9018 12070 9110 12162
<< locali >>
rect 1709 23198 1735 23243
rect 441 20345 442 20407
rect 1709 19934 1735 19979
rect 441 17081 442 17143
rect 1709 16670 1735 16715
rect 441 13817 442 13879
rect 1709 13406 1735 13451
rect 9693 11687 9746 11811
rect 11631 11701 11665 11746
rect 441 10553 442 10615
rect 1709 10142 1735 10187
rect 441 7289 442 7351
rect 1709 6878 1735 6923
rect 441 4025 442 4087
<< viali >>
rect 1769 23209 1803 23243
rect 442 20345 504 20407
rect 1769 19945 1803 19979
rect 442 17081 504 17143
rect 1769 16681 1803 16715
rect 442 13817 504 13879
rect 1769 13417 1803 13451
rect 9071 11637 9137 11703
rect 9257 11678 9325 11746
rect 9442 11684 9498 11740
rect 9890 11737 9964 11811
rect 10369 11741 10429 11801
rect 10676 11749 10725 11798
rect 10927 11737 10985 11795
rect 442 10553 504 10615
rect 1769 10153 1803 10187
rect 442 7289 504 7351
rect 1769 6889 1803 6923
rect 442 4025 504 4087
rect 1769 3625 1803 3659
rect 442 761 504 823
<< metal1 >>
rect 1763 23243 1815 23249
rect 438 23184 444 23243
rect 503 23209 1769 23243
rect 1803 23209 1815 23243
rect 503 23184 509 23209
rect 1763 23203 1815 23209
rect 436 20413 510 20419
rect 430 20351 436 20413
rect 510 20351 516 20413
rect 430 20345 442 20351
rect 504 20345 516 20351
rect 430 20339 516 20345
rect 1763 19979 1815 19985
rect 438 19920 444 19979
rect 503 19945 1769 19979
rect 1803 19945 1815 19979
rect 503 19920 509 19945
rect 1763 19939 1815 19945
rect 436 17149 510 17155
rect 430 17087 436 17149
rect 510 17087 516 17149
rect 430 17081 442 17087
rect 504 17081 516 17087
rect 430 17075 516 17081
rect 1763 16715 1815 16721
rect 438 16656 444 16715
rect 503 16681 1769 16715
rect 1803 16681 1815 16715
rect 503 16656 509 16681
rect 1763 16675 1815 16681
rect 436 13885 510 13891
rect 430 13823 436 13885
rect 510 13823 516 13885
rect 430 13817 442 13823
rect 504 13817 516 13823
rect 430 13811 516 13817
rect 1763 13451 1815 13457
rect 438 13392 444 13451
rect 503 13417 1769 13451
rect 1803 13417 1815 13451
rect 503 13392 509 13417
rect 1763 13411 1815 13417
rect 9884 11811 9970 11823
rect 9884 11805 9890 11811
rect 9964 11805 9970 11811
rect 8950 11612 8956 11790
rect 9134 11709 9140 11790
rect 9245 11746 9331 11752
rect 9134 11703 9143 11709
rect 9137 11637 9143 11703
rect 9245 11678 9257 11746
rect 9325 11740 9510 11746
rect 9325 11684 9442 11740
rect 9498 11684 9510 11740
rect 10357 11801 10441 11807
rect 10357 11795 10369 11801
rect 10429 11795 10441 11801
rect 10357 11735 10363 11795
rect 10435 11735 10441 11795
rect 10664 11798 10737 11804
rect 10664 11795 10676 11798
rect 10725 11795 10737 11798
rect 10664 11743 10670 11795
rect 10731 11743 10737 11795
rect 10670 11737 10731 11743
rect 9884 11725 9970 11731
rect 10363 11729 10435 11735
rect 10915 11731 10921 11801
rect 10991 11731 10997 11801
rect 9325 11678 9510 11684
rect 9245 11677 9331 11678
rect 9251 11672 9331 11677
rect 9134 11631 9143 11637
rect 9134 11612 9140 11631
rect 436 10621 510 10627
rect 430 10559 436 10621
rect 510 10559 516 10621
rect 430 10553 442 10559
rect 504 10553 516 10559
rect 430 10547 516 10553
rect 1763 10187 1815 10193
rect 438 10128 444 10187
rect 503 10153 1769 10187
rect 1803 10153 1815 10187
rect 503 10128 509 10153
rect 1763 10147 1815 10153
rect 436 7357 510 7363
rect 430 7295 436 7357
rect 510 7295 516 7357
rect 430 7289 442 7295
rect 504 7289 516 7295
rect 430 7283 516 7289
rect 1763 6923 1815 6929
rect 438 6864 444 6923
rect 503 6889 1769 6923
rect 1803 6889 1815 6923
rect 503 6864 509 6889
rect 1763 6883 1815 6889
rect 436 4093 510 4099
rect 430 4031 436 4093
rect 510 4031 516 4093
rect 430 4025 442 4031
rect 504 4025 516 4031
rect 430 4019 516 4025
rect 1763 3659 1815 3665
rect 438 3600 444 3659
rect 503 3625 1769 3659
rect 1803 3625 1815 3659
rect 503 3600 509 3625
rect 1763 3619 1815 3625
rect 436 829 510 835
rect 430 767 436 829
rect 510 767 516 829
rect 430 761 442 767
rect 504 761 516 767
rect 430 755 516 761
<< via1 >>
rect 444 23184 503 23243
rect 436 20407 510 20413
rect 436 20351 442 20407
rect 442 20351 504 20407
rect 504 20351 510 20407
rect 444 19920 503 19979
rect 436 17143 510 17149
rect 436 17087 442 17143
rect 442 17087 504 17143
rect 504 17087 510 17143
rect 444 16656 503 16715
rect 436 13879 510 13885
rect 436 13823 442 13879
rect 442 13823 504 13879
rect 504 13823 510 13879
rect 444 13392 503 13451
rect 8956 11703 9134 11790
rect 8956 11637 9071 11703
rect 9071 11637 9134 11703
rect 9884 11737 9890 11805
rect 9890 11737 9964 11805
rect 9964 11737 9970 11805
rect 9884 11731 9970 11737
rect 10363 11741 10369 11795
rect 10369 11741 10429 11795
rect 10429 11741 10435 11795
rect 10363 11735 10435 11741
rect 10670 11749 10676 11795
rect 10676 11749 10725 11795
rect 10725 11749 10731 11795
rect 10670 11743 10731 11749
rect 10921 11795 10991 11801
rect 10921 11737 10927 11795
rect 10927 11737 10985 11795
rect 10985 11737 10991 11795
rect 10921 11731 10991 11737
rect 8956 11612 9134 11637
rect 436 10615 510 10621
rect 436 10559 442 10615
rect 442 10559 504 10615
rect 504 10559 510 10615
rect 444 10128 503 10187
rect 436 7351 510 7357
rect 436 7295 442 7351
rect 442 7295 504 7351
rect 504 7295 510 7351
rect 444 6864 503 6923
rect 436 4087 510 4093
rect 436 4031 442 4087
rect 442 4031 504 4087
rect 504 4031 510 4087
rect 444 3600 503 3659
rect 436 823 510 829
rect 436 767 442 823
rect 442 767 504 823
rect 504 767 510 823
<< metal2 >>
rect 444 23243 503 23249
rect 444 20413 503 23184
rect 6046 22935 6142 23504
rect -276 20351 436 20413
rect 510 20351 516 20413
rect -276 16 -217 20351
rect 444 20339 503 20351
rect 444 19979 503 19985
rect 444 17149 503 19920
rect -156 17087 436 17149
rect 510 17087 516 17149
rect -156 16 -97 17087
rect 444 17075 503 17087
rect 444 16715 503 16721
rect 444 13885 503 16656
rect -36 13823 436 13885
rect 510 13823 516 13885
rect -36 16 23 13823
rect 444 13811 503 13823
rect 444 13451 503 13457
rect 444 10621 503 13392
rect 8956 11790 9134 11796
rect 6001 11612 8529 11790
rect 8707 11612 8716 11790
rect 9878 11731 9884 11805
rect 9970 11731 9976 11805
rect 10921 11801 10991 11807
rect 10357 11735 10363 11795
rect 10435 11735 10441 11795
rect 10664 11743 10670 11795
rect 10731 11743 10737 11795
rect 8956 11606 9134 11612
rect 9890 11440 9964 11731
rect 10369 11440 10429 11735
rect 10676 11440 10725 11743
rect 10921 11725 10991 11731
rect 10927 11440 10985 11725
rect 84 10559 436 10621
rect 510 10559 516 10621
rect 84 16 143 10559
rect 444 10547 503 10559
rect 444 10187 503 10193
rect 444 7357 503 10128
rect 204 7295 436 7357
rect 510 7295 516 7357
rect 204 16 263 7295
rect 444 7283 503 7295
rect 444 6923 503 6929
rect 444 4093 503 6864
rect 324 4031 436 4093
rect 510 4031 516 4093
rect 324 16 383 4031
rect 444 4019 503 4031
rect 444 3659 503 3665
rect 444 829 503 3600
rect 430 767 436 829
rect 510 767 516 829
rect 444 16 503 767
<< via2 >>
rect 8529 11612 8707 11790
rect 8961 11617 9129 11785
<< metal3 >>
rect 8524 11790 8712 11795
rect 8524 11612 8529 11790
rect 8707 11785 9134 11790
rect 8707 11617 8961 11785
rect 9129 11617 9134 11785
rect 8707 11612 9134 11617
rect 8524 11607 8712 11612
use SSTL  SSTL_0 ~/proj/caravan-project/mag/SSTL
timestamp 1644115763
transform 1 0 2350 0 -1 4308
box -2332 -19196 6668 4292
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 8980 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_1
timestamp 1644111581
transform 1 0 9348 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 11648 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 9716 0 1 11488
box -38 -48 1970 592
<< end >>
