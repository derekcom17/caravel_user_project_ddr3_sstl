magic
tech sky130A
magscale 1 2
timestamp 1644853372
<< nwell >>
rect 20242 32742 20626 32834
rect 20242 29478 20626 29570
rect 20242 26214 20626 26306
rect 20242 22950 20626 23042
rect 20242 19686 20626 19778
rect 20242 16422 20626 16514
rect 20242 13158 20626 13250
rect 9018 12070 9110 12162
<< locali >>
rect 19819 32313 20159 32425
rect 19819 29049 20159 29161
rect 19819 25785 20159 25897
rect 1709 23198 1735 23243
rect 19819 22521 20159 22633
rect 441 20345 442 20407
rect 1709 19934 1735 19979
rect 19819 19257 20159 19369
rect 441 17081 442 17143
rect 1709 16670 1735 16715
rect 19819 15993 20159 16105
rect 441 13817 442 13879
rect 1709 13406 1735 13451
rect 19819 12729 20159 12841
rect 9693 11687 9746 11811
rect 11631 11701 11665 11746
rect 441 10553 442 10615
rect 1709 10142 1735 10187
rect 441 7289 442 7351
rect 1709 6878 1735 6923
rect 441 4025 442 4087
<< viali >>
rect 18463 35167 18501 35205
rect 20221 35161 20271 35211
rect 22377 35166 22411 35200
rect 20159 32313 20271 32425
rect 21062 32314 21106 32358
rect 18463 31903 18501 31941
rect 20221 31897 20271 31947
rect 22377 31902 22411 31936
rect 20159 29049 20271 29161
rect 21062 29050 21106 29094
rect 18463 28639 18501 28677
rect 20221 28633 20271 28683
rect 22377 28638 22411 28672
rect 20159 25785 20271 25897
rect 21062 25786 21106 25830
rect 18463 25375 18501 25413
rect 20221 25369 20271 25419
rect 22377 25374 22411 25408
rect 1769 23209 1803 23243
rect 20159 22521 20271 22633
rect 21062 22522 21106 22566
rect 18463 22111 18501 22149
rect 20221 22105 20271 22155
rect 22377 22110 22411 22144
rect 442 20345 504 20407
rect 1769 19945 1803 19979
rect 20159 19257 20271 19369
rect 21062 19258 21106 19302
rect 18463 18847 18501 18885
rect 20221 18841 20271 18891
rect 22377 18846 22411 18880
rect 442 17081 504 17143
rect 1769 16681 1803 16715
rect 20159 15993 20271 16105
rect 21062 15994 21106 16038
rect 18463 15583 18501 15621
rect 20221 15577 20271 15627
rect 22377 15582 22411 15616
rect 442 13817 504 13879
rect 1769 13417 1803 13451
rect 20159 12729 20271 12841
rect 21062 12730 21106 12774
rect 9071 11637 9137 11703
rect 9257 11678 9325 11746
rect 9442 11684 9498 11740
rect 9890 11737 9964 11811
rect 10369 11741 10429 11801
rect 10676 11749 10725 11798
rect 10927 11737 10985 11795
rect 442 10553 504 10615
rect 1769 10153 1803 10187
rect 442 7289 504 7351
rect 1769 6889 1803 6923
rect 442 4025 504 4087
rect 1769 3625 1803 3659
rect 442 761 504 823
<< metal1 >>
rect 20215 35211 20277 35223
rect 18451 35205 20221 35211
rect 18451 35167 18463 35205
rect 18501 35167 20221 35205
rect 18451 35161 20221 35167
rect 20271 35183 20277 35211
rect 20908 35183 20964 35189
rect 20271 35161 20908 35183
rect 20215 35149 20908 35161
rect 20221 35127 20908 35149
rect 21001 35140 21007 35253
rect 21120 35209 21126 35253
rect 21124 35200 21130 35209
rect 22365 35200 22423 35206
rect 21124 35166 22377 35200
rect 22411 35166 22423 35200
rect 21124 35157 21130 35166
rect 22365 35160 22423 35166
rect 21120 35140 21126 35157
rect 20908 35121 20964 35127
rect 21007 32585 21120 32591
rect 20159 32472 21007 32585
rect 20159 32437 20272 32472
rect 21007 32466 21120 32472
rect 20153 32425 20277 32437
rect 20153 32313 20159 32425
rect 20271 32313 20277 32425
rect 20153 32301 20277 32313
rect 20902 32308 20908 32364
rect 20964 32358 21118 32364
rect 20964 32314 21062 32358
rect 21106 32314 21118 32358
rect 20964 32308 21118 32314
rect 20215 31947 20277 31959
rect 18451 31941 20221 31947
rect 18451 31903 18463 31941
rect 18501 31903 20221 31941
rect 18451 31897 20221 31903
rect 20271 31919 20277 31947
rect 20908 31919 20964 31925
rect 20271 31897 20908 31919
rect 20215 31885 20908 31897
rect 20221 31863 20908 31885
rect 21001 31876 21007 31989
rect 21120 31945 21126 31989
rect 21124 31936 21130 31945
rect 22365 31936 22423 31942
rect 21124 31902 22377 31936
rect 22411 31902 22423 31936
rect 21124 31893 21130 31902
rect 22365 31896 22423 31902
rect 21120 31876 21126 31893
rect 20908 31857 20964 31863
rect 21007 29321 21120 29327
rect 20159 29208 21007 29321
rect 20159 29173 20272 29208
rect 21007 29202 21120 29208
rect 20153 29161 20277 29173
rect 20153 29049 20159 29161
rect 20271 29049 20277 29161
rect 20153 29037 20277 29049
rect 20902 29044 20908 29100
rect 20964 29094 21118 29100
rect 20964 29050 21062 29094
rect 21106 29050 21118 29094
rect 20964 29044 21118 29050
rect 20215 28683 20277 28695
rect 18451 28677 20221 28683
rect 18451 28639 18463 28677
rect 18501 28639 20221 28677
rect 18451 28633 20221 28639
rect 20271 28655 20277 28683
rect 20908 28655 20964 28661
rect 20271 28633 20908 28655
rect 20215 28621 20908 28633
rect 20221 28599 20908 28621
rect 21001 28612 21007 28725
rect 21120 28681 21126 28725
rect 21124 28672 21130 28681
rect 22365 28672 22423 28678
rect 21124 28638 22377 28672
rect 22411 28638 22423 28672
rect 21124 28629 21130 28638
rect 22365 28632 22423 28638
rect 21120 28612 21126 28629
rect 20908 28593 20964 28599
rect 21007 26057 21120 26063
rect 20159 25944 21007 26057
rect 20159 25909 20272 25944
rect 21007 25938 21120 25944
rect 20153 25897 20277 25909
rect 20153 25785 20159 25897
rect 20271 25785 20277 25897
rect 20153 25773 20277 25785
rect 20902 25780 20908 25836
rect 20964 25830 21118 25836
rect 20964 25786 21062 25830
rect 21106 25786 21118 25830
rect 20964 25780 21118 25786
rect 20215 25419 20277 25431
rect 18451 25413 20221 25419
rect 18451 25375 18463 25413
rect 18501 25375 20221 25413
rect 18451 25369 20221 25375
rect 20271 25391 20277 25419
rect 20908 25391 20964 25397
rect 20271 25369 20908 25391
rect 20215 25357 20908 25369
rect 20221 25335 20908 25357
rect 21001 25348 21007 25461
rect 21120 25417 21126 25461
rect 21124 25408 21130 25417
rect 22365 25408 22423 25414
rect 21124 25374 22377 25408
rect 22411 25374 22423 25408
rect 21124 25365 21130 25374
rect 22365 25368 22423 25374
rect 21120 25348 21126 25365
rect 20908 25329 20964 25335
rect 1763 23243 1815 23249
rect 438 23184 444 23243
rect 503 23209 1769 23243
rect 1803 23209 1815 23243
rect 503 23184 509 23209
rect 1763 23203 1815 23209
rect 21007 22793 21120 22799
rect 20159 22680 21007 22793
rect 20159 22645 20272 22680
rect 21007 22674 21120 22680
rect 20153 22633 20277 22645
rect 20153 22521 20159 22633
rect 20271 22521 20277 22633
rect 20153 22509 20277 22521
rect 20902 22516 20908 22572
rect 20964 22566 21118 22572
rect 20964 22522 21062 22566
rect 21106 22522 21118 22566
rect 20964 22516 21118 22522
rect 20215 22155 20277 22167
rect 18451 22149 20221 22155
rect 18451 22111 18463 22149
rect 18501 22111 20221 22149
rect 18451 22105 20221 22111
rect 20271 22127 20277 22155
rect 20908 22127 20964 22133
rect 20271 22105 20908 22127
rect 20215 22093 20908 22105
rect 20221 22071 20908 22093
rect 21001 22084 21007 22197
rect 21120 22153 21126 22197
rect 21124 22144 21130 22153
rect 22365 22144 22423 22150
rect 21124 22110 22377 22144
rect 22411 22110 22423 22144
rect 21124 22101 21130 22110
rect 22365 22104 22423 22110
rect 21120 22084 21126 22101
rect 20908 22065 20964 22071
rect 436 20413 510 20419
rect 430 20351 436 20413
rect 510 20351 516 20413
rect 430 20345 442 20351
rect 504 20345 516 20351
rect 430 20339 516 20345
rect 1763 19979 1815 19985
rect 438 19920 444 19979
rect 503 19945 1769 19979
rect 1803 19945 1815 19979
rect 503 19920 509 19945
rect 1763 19939 1815 19945
rect 21007 19529 21120 19535
rect 20159 19416 21007 19529
rect 20159 19381 20272 19416
rect 21007 19410 21120 19416
rect 20153 19369 20277 19381
rect 20153 19257 20159 19369
rect 20271 19257 20277 19369
rect 20153 19245 20277 19257
rect 20902 19252 20908 19308
rect 20964 19302 21118 19308
rect 20964 19258 21062 19302
rect 21106 19258 21118 19302
rect 20964 19252 21118 19258
rect 20215 18891 20277 18903
rect 18451 18885 20221 18891
rect 18451 18847 18463 18885
rect 18501 18847 20221 18885
rect 18451 18841 20221 18847
rect 20271 18863 20277 18891
rect 20908 18863 20964 18869
rect 20271 18841 20908 18863
rect 20215 18829 20908 18841
rect 20221 18807 20908 18829
rect 21001 18820 21007 18933
rect 21120 18889 21126 18933
rect 21124 18880 21130 18889
rect 22365 18880 22423 18886
rect 21124 18846 22377 18880
rect 22411 18846 22423 18880
rect 21124 18837 21130 18846
rect 22365 18840 22423 18846
rect 21120 18820 21126 18837
rect 20908 18801 20964 18807
rect 436 17149 510 17155
rect 430 17087 436 17149
rect 510 17087 516 17149
rect 430 17081 442 17087
rect 504 17081 516 17087
rect 430 17075 516 17081
rect 1763 16715 1815 16721
rect 438 16656 444 16715
rect 503 16681 1769 16715
rect 1803 16681 1815 16715
rect 503 16656 509 16681
rect 1763 16675 1815 16681
rect 21007 16265 21120 16271
rect 20159 16152 21007 16265
rect 20159 16117 20272 16152
rect 21007 16146 21120 16152
rect 20153 16105 20277 16117
rect 20153 15993 20159 16105
rect 20271 15993 20277 16105
rect 20153 15981 20277 15993
rect 20902 15988 20908 16044
rect 20964 16038 21118 16044
rect 20964 15994 21062 16038
rect 21106 15994 21118 16038
rect 20964 15988 21118 15994
rect 20215 15627 20277 15639
rect 18451 15621 20221 15627
rect 18451 15583 18463 15621
rect 18501 15583 20221 15621
rect 18451 15577 20221 15583
rect 20271 15599 20277 15627
rect 20908 15599 20964 15605
rect 20271 15577 20908 15599
rect 20215 15565 20908 15577
rect 20221 15543 20908 15565
rect 21001 15556 21007 15669
rect 21120 15625 21126 15669
rect 21124 15616 21130 15625
rect 22365 15616 22423 15622
rect 21124 15582 22377 15616
rect 22411 15582 22423 15616
rect 21124 15573 21130 15582
rect 22365 15576 22423 15582
rect 21120 15556 21126 15573
rect 20908 15537 20964 15543
rect 436 13885 510 13891
rect 430 13823 436 13885
rect 510 13823 516 13885
rect 430 13817 442 13823
rect 504 13817 516 13823
rect 430 13811 516 13817
rect 1763 13451 1815 13457
rect 438 13392 444 13451
rect 503 13417 1769 13451
rect 1803 13417 1815 13451
rect 503 13392 509 13417
rect 1763 13411 1815 13417
rect 21007 13001 21120 13007
rect 20159 12888 21007 13001
rect 20159 12853 20272 12888
rect 21007 12882 21120 12888
rect 20153 12841 20277 12853
rect 20153 12729 20159 12841
rect 20271 12729 20277 12841
rect 20153 12717 20277 12729
rect 20902 12724 20908 12780
rect 20964 12774 21118 12780
rect 20964 12730 21062 12774
rect 21106 12730 21118 12774
rect 20964 12724 21118 12730
rect 9884 11811 9970 11823
rect 9884 11805 9890 11811
rect 9964 11805 9970 11811
rect 9245 11746 9331 11752
rect 6024 11617 6030 11724
rect 6137 11703 9158 11724
rect 6137 11637 9071 11703
rect 9137 11637 9158 11703
rect 9245 11678 9257 11746
rect 9325 11740 9510 11746
rect 9325 11684 9442 11740
rect 9498 11684 9510 11740
rect 10357 11801 10441 11807
rect 10357 11795 10369 11801
rect 10429 11795 10441 11801
rect 10357 11735 10363 11795
rect 10435 11735 10441 11795
rect 10664 11798 10737 11804
rect 10664 11795 10676 11798
rect 10725 11795 10737 11798
rect 10664 11743 10670 11795
rect 10731 11743 10737 11795
rect 10670 11737 10731 11743
rect 9884 11725 9970 11731
rect 10363 11729 10435 11735
rect 10915 11731 10921 11801
rect 10991 11731 10997 11801
rect 9325 11678 9510 11684
rect 9245 11677 9331 11678
rect 9251 11672 9331 11677
rect 6137 11617 9158 11637
rect 436 10621 510 10627
rect 430 10559 436 10621
rect 510 10559 516 10621
rect 430 10553 442 10559
rect 504 10553 516 10559
rect 430 10547 516 10553
rect 1763 10187 1815 10193
rect 438 10128 444 10187
rect 503 10153 1769 10187
rect 1803 10153 1815 10187
rect 503 10128 509 10153
rect 1763 10147 1815 10153
rect 436 7357 510 7363
rect 430 7295 436 7357
rect 510 7295 516 7357
rect 430 7289 442 7295
rect 504 7289 516 7295
rect 430 7283 516 7289
rect 1763 6923 1815 6929
rect 438 6864 444 6923
rect 503 6889 1769 6923
rect 1803 6889 1815 6923
rect 503 6864 509 6889
rect 1763 6883 1815 6889
rect 436 4093 510 4099
rect 430 4031 436 4093
rect 510 4031 516 4093
rect 430 4025 442 4031
rect 504 4025 516 4031
rect 430 4019 516 4025
rect 1763 3659 1815 3665
rect 438 3600 444 3659
rect 503 3625 1769 3659
rect 1803 3625 1815 3659
rect 503 3600 509 3625
rect 1763 3619 1815 3625
rect 436 829 510 835
rect 430 767 436 829
rect 510 767 516 829
rect 430 761 442 767
rect 504 761 516 767
rect 430 755 516 761
<< via1 >>
rect 20908 35127 20964 35183
rect 21007 35209 21120 35253
rect 21007 35157 21124 35209
rect 21007 35140 21120 35157
rect 21007 32472 21120 32585
rect 20908 32308 20964 32364
rect 20908 31863 20964 31919
rect 21007 31945 21120 31989
rect 21007 31893 21124 31945
rect 21007 31876 21120 31893
rect 21007 29208 21120 29321
rect 20908 29044 20964 29100
rect 20908 28599 20964 28655
rect 21007 28681 21120 28725
rect 21007 28629 21124 28681
rect 21007 28612 21120 28629
rect 21007 25944 21120 26057
rect 20908 25780 20964 25836
rect 20908 25335 20964 25391
rect 21007 25417 21120 25461
rect 21007 25365 21124 25417
rect 21007 25348 21120 25365
rect 444 23184 503 23243
rect 21007 22680 21120 22793
rect 20908 22516 20964 22572
rect 20908 22071 20964 22127
rect 21007 22153 21120 22197
rect 21007 22101 21124 22153
rect 21007 22084 21120 22101
rect 436 20407 510 20413
rect 436 20351 442 20407
rect 442 20351 504 20407
rect 504 20351 510 20407
rect 444 19920 503 19979
rect 21007 19416 21120 19529
rect 20908 19252 20964 19308
rect 20908 18807 20964 18863
rect 21007 18889 21120 18933
rect 21007 18837 21124 18889
rect 21007 18820 21120 18837
rect 436 17143 510 17149
rect 436 17087 442 17143
rect 442 17087 504 17143
rect 504 17087 510 17143
rect 444 16656 503 16715
rect 21007 16152 21120 16265
rect 20908 15988 20964 16044
rect 20908 15543 20964 15599
rect 21007 15625 21120 15669
rect 21007 15573 21124 15625
rect 21007 15556 21120 15573
rect 436 13879 510 13885
rect 436 13823 442 13879
rect 442 13823 504 13879
rect 504 13823 510 13879
rect 444 13392 503 13451
rect 21007 12888 21120 13001
rect 20908 12724 20964 12780
rect 6030 11617 6137 11724
rect 9884 11737 9890 11805
rect 9890 11737 9964 11805
rect 9964 11737 9970 11805
rect 9884 11731 9970 11737
rect 10363 11741 10369 11795
rect 10369 11741 10429 11795
rect 10429 11741 10435 11795
rect 10363 11735 10435 11741
rect 10670 11749 10676 11795
rect 10676 11749 10725 11795
rect 10725 11749 10731 11795
rect 10670 11743 10731 11749
rect 10921 11795 10991 11801
rect 10921 11737 10927 11795
rect 10927 11737 10985 11795
rect 10985 11737 10991 11795
rect 10921 11731 10991 11737
rect 436 10615 510 10621
rect 436 10559 442 10615
rect 442 10559 504 10615
rect 504 10559 510 10615
rect 444 10128 503 10187
rect 436 7351 510 7357
rect 436 7295 442 7351
rect 442 7295 504 7351
rect 504 7295 510 7351
rect 444 6864 503 6923
rect 436 4087 510 4093
rect 436 4031 442 4087
rect 442 4031 504 4087
rect 504 4031 510 4087
rect 444 3600 503 3659
rect 436 823 510 829
rect 436 767 442 823
rect 442 767 504 823
rect 504 767 510 823
<< metal2 >>
rect 21007 35253 21120 35259
rect 21120 35209 21124 35215
rect 20902 35127 20908 35183
rect 20964 35127 20970 35183
rect 21120 35151 21124 35157
rect 20908 32364 20964 35127
rect 21007 32585 21120 35140
rect 21001 32472 21007 32585
rect 21120 32472 21126 32585
rect 20908 32302 20964 32308
rect 21007 31989 21120 31995
rect 21120 31945 21124 31951
rect 20902 31863 20908 31919
rect 20964 31863 20970 31919
rect 21120 31887 21124 31893
rect 20908 29100 20964 31863
rect 21007 29321 21120 31876
rect 21001 29208 21007 29321
rect 21120 29208 21126 29321
rect 20908 29038 20964 29044
rect 21007 28725 21120 28731
rect 21120 28681 21124 28687
rect 20902 28599 20908 28655
rect 20964 28599 20970 28655
rect 21120 28623 21124 28629
rect 20908 25836 20964 28599
rect 21007 26057 21120 28612
rect 21001 25944 21007 26057
rect 21120 25944 21126 26057
rect 20908 25774 20964 25780
rect 21007 25461 21120 25467
rect 21120 25417 21124 25423
rect 20902 25335 20908 25391
rect 20964 25335 20970 25391
rect 21120 25359 21124 25365
rect 444 23243 503 23249
rect 444 20413 503 23184
rect 6046 22935 6142 23504
rect 20908 22572 20964 25335
rect 21007 22793 21120 25348
rect 21001 22680 21007 22793
rect 21120 22680 21126 22793
rect 20908 22510 20964 22516
rect 21007 22197 21120 22203
rect 21120 22153 21124 22159
rect 20902 22071 20908 22127
rect 20964 22071 20970 22127
rect 21120 22095 21124 22101
rect -276 20351 436 20413
rect 510 20351 516 20413
rect -276 16 -217 20351
rect 444 20339 503 20351
rect 444 19979 503 19985
rect 444 17149 503 19920
rect 20908 19308 20964 22071
rect 21007 19529 21120 22084
rect 21001 19416 21007 19529
rect 21120 19416 21126 19529
rect 20908 19246 20964 19252
rect 21007 18933 21120 18939
rect 21120 18889 21124 18895
rect 20902 18807 20908 18863
rect 20964 18807 20970 18863
rect 21120 18831 21124 18837
rect -156 17087 436 17149
rect 510 17087 516 17149
rect -156 16 -97 17087
rect 444 17075 503 17087
rect 444 16715 503 16721
rect 444 13885 503 16656
rect 20908 16044 20964 18807
rect 21007 16265 21120 18820
rect 21001 16152 21007 16265
rect 21120 16152 21126 16265
rect 20908 15982 20964 15988
rect 21007 15669 21120 15675
rect 21120 15625 21124 15631
rect 20902 15543 20908 15599
rect 20964 15543 20970 15599
rect 21120 15567 21124 15573
rect -36 13823 436 13885
rect 510 13823 516 13885
rect -36 16 23 13823
rect 444 13811 503 13823
rect 444 13451 503 13457
rect 444 10621 503 13392
rect 20908 12780 20964 15543
rect 21007 13001 21120 15556
rect 21001 12888 21007 13001
rect 21120 12888 21126 13001
rect 20908 12718 20964 12724
rect 9878 11731 9884 11805
rect 9970 11731 9976 11805
rect 10921 11801 10991 11807
rect 10357 11735 10363 11795
rect 10435 11735 10441 11795
rect 10664 11743 10670 11795
rect 10731 11743 10737 11795
rect 6030 11724 6137 11730
rect 6030 11611 6137 11617
rect 9890 11440 9964 11731
rect 10369 11440 10429 11735
rect 10676 11440 10725 11743
rect 10921 11725 10991 11731
rect 10927 11440 10985 11725
rect 84 10559 436 10621
rect 510 10559 516 10621
rect 84 16 143 10559
rect 444 10547 503 10559
rect 444 10187 503 10193
rect 444 7357 503 10128
rect 204 7295 436 7357
rect 510 7295 516 7357
rect 204 16 263 7295
rect 444 7283 503 7295
rect 444 6923 503 6929
rect 444 4093 503 6864
rect 324 4031 436 4093
rect 510 4031 516 4093
rect 324 16 383 4031
rect 444 4019 503 4031
rect 444 3659 503 3665
rect 444 829 503 3600
rect 430 767 436 829
rect 510 767 516 829
rect 444 16 503 767
use SSTL  SSTL_0 ~/proj/caravan-project/mag/SSTL
timestamp 1644115763
transform 1 0 2350 0 -1 4308
box -2332 -19196 6668 4292
use SSTL  SSTL_1
timestamp 1644115763
transform -1 0 17910 0 -1 16276
box -2332 -19196 6668 4292
use SSTL  SSTL_2
timestamp 1644115763
transform 1 0 22958 0 -1 16276
box -2332 -19196 6668 4292
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform -1 0 20664 0 1 12576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1644111581
transform -1 0 20664 0 -1 15840
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1644111581
transform -1 0 20664 0 -1 19104
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1644111581
transform -1 0 20664 0 1 15840
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1644111581
transform -1 0 20664 0 -1 22368
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1644111581
transform -1 0 20664 0 1 19104
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1644111581
transform -1 0 20664 0 -1 25632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_7
timestamp 1644111581
transform -1 0 20664 0 1 22368
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_8
timestamp 1644111581
transform -1 0 20664 0 -1 28896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_9
timestamp 1644111581
transform -1 0 20664 0 1 25632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_10
timestamp 1644111581
transform -1 0 20664 0 -1 32160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_11
timestamp 1644111581
transform -1 0 20664 0 1 28896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_12
timestamp 1644111581
transform -1 0 20664 0 -1 35424
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_13
timestamp 1644111581
transform -1 0 20664 0 1 32160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 8980 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_1
timestamp 1644111581
transform 1 0 9348 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 11648 0 1 11488
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 ~/proj/caravan-project/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644111581
transform 1 0 9716 0 1 11488
box -38 -48 1970 592
<< end >>
